library ieee;
use ieee.std_logic_1164.all;

package types is
    -- FUNCTIONS

    -- CONSTANTS

    -- DATA TYPES
    type bus_array is array(15 downto 0) of signed (7 downto 0);

end package;


-- FUNCTION DEFINITIONS
-- package body types is
    
--     function x (a:integer, b:integer) return integer is
--     begin
--         ...
--     end x;

-- end package body;
