-- dma_platform.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity dma_platform is
	port (
		arm_a9_hps_f2h_stm_hw_events_stm_hwevents : in    std_logic_vector(27 downto 0) := (others => '0'); -- arm_a9_hps_f2h_stm_hw_events.stm_hwevents
		hps_io_hps_io_emac1_inst_TX_CLK           : out   std_logic;                                        --                       hps_io.hps_io_emac1_inst_TX_CLK
		hps_io_hps_io_emac1_inst_TXD0             : out   std_logic;                                        --                             .hps_io_emac1_inst_TXD0
		hps_io_hps_io_emac1_inst_TXD1             : out   std_logic;                                        --                             .hps_io_emac1_inst_TXD1
		hps_io_hps_io_emac1_inst_TXD2             : out   std_logic;                                        --                             .hps_io_emac1_inst_TXD2
		hps_io_hps_io_emac1_inst_TXD3             : out   std_logic;                                        --                             .hps_io_emac1_inst_TXD3
		hps_io_hps_io_emac1_inst_RXD0             : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RXD0
		hps_io_hps_io_emac1_inst_MDIO             : inout std_logic                     := '0';             --                             .hps_io_emac1_inst_MDIO
		hps_io_hps_io_emac1_inst_MDC              : out   std_logic;                                        --                             .hps_io_emac1_inst_MDC
		hps_io_hps_io_emac1_inst_RX_CTL           : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RX_CTL
		hps_io_hps_io_emac1_inst_TX_CTL           : out   std_logic;                                        --                             .hps_io_emac1_inst_TX_CTL
		hps_io_hps_io_emac1_inst_RX_CLK           : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RX_CLK
		hps_io_hps_io_emac1_inst_RXD1             : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RXD1
		hps_io_hps_io_emac1_inst_RXD2             : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RXD2
		hps_io_hps_io_emac1_inst_RXD3             : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RXD3
		hps_io_hps_io_qspi_inst_IO0               : inout std_logic                     := '0';             --                             .hps_io_qspi_inst_IO0
		hps_io_hps_io_qspi_inst_IO1               : inout std_logic                     := '0';             --                             .hps_io_qspi_inst_IO1
		hps_io_hps_io_qspi_inst_IO2               : inout std_logic                     := '0';             --                             .hps_io_qspi_inst_IO2
		hps_io_hps_io_qspi_inst_IO3               : inout std_logic                     := '0';             --                             .hps_io_qspi_inst_IO3
		hps_io_hps_io_qspi_inst_SS0               : out   std_logic;                                        --                             .hps_io_qspi_inst_SS0
		hps_io_hps_io_qspi_inst_CLK               : out   std_logic;                                        --                             .hps_io_qspi_inst_CLK
		hps_io_hps_io_sdio_inst_CMD               : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_CMD
		hps_io_hps_io_sdio_inst_D0                : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_D0
		hps_io_hps_io_sdio_inst_D1                : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_D1
		hps_io_hps_io_sdio_inst_CLK               : out   std_logic;                                        --                             .hps_io_sdio_inst_CLK
		hps_io_hps_io_sdio_inst_D2                : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_D2
		hps_io_hps_io_sdio_inst_D3                : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_D3
		hps_io_hps_io_usb1_inst_D0                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D0
		hps_io_hps_io_usb1_inst_D1                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D1
		hps_io_hps_io_usb1_inst_D2                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D2
		hps_io_hps_io_usb1_inst_D3                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D3
		hps_io_hps_io_usb1_inst_D4                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D4
		hps_io_hps_io_usb1_inst_D5                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D5
		hps_io_hps_io_usb1_inst_D6                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D6
		hps_io_hps_io_usb1_inst_D7                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D7
		hps_io_hps_io_usb1_inst_CLK               : in    std_logic                     := '0';             --                             .hps_io_usb1_inst_CLK
		hps_io_hps_io_usb1_inst_STP               : out   std_logic;                                        --                             .hps_io_usb1_inst_STP
		hps_io_hps_io_usb1_inst_DIR               : in    std_logic                     := '0';             --                             .hps_io_usb1_inst_DIR
		hps_io_hps_io_usb1_inst_NXT               : in    std_logic                     := '0';             --                             .hps_io_usb1_inst_NXT
		hps_io_hps_io_spim0_inst_CLK              : out   std_logic;                                        --                             .hps_io_spim0_inst_CLK
		hps_io_hps_io_spim0_inst_MOSI             : out   std_logic;                                        --                             .hps_io_spim0_inst_MOSI
		hps_io_hps_io_spim0_inst_MISO             : in    std_logic                     := '0';             --                             .hps_io_spim0_inst_MISO
		hps_io_hps_io_spim0_inst_SS0              : out   std_logic;                                        --                             .hps_io_spim0_inst_SS0
		hps_io_hps_io_spim1_inst_CLK              : out   std_logic;                                        --                             .hps_io_spim1_inst_CLK
		hps_io_hps_io_spim1_inst_MOSI             : out   std_logic;                                        --                             .hps_io_spim1_inst_MOSI
		hps_io_hps_io_spim1_inst_MISO             : in    std_logic                     := '0';             --                             .hps_io_spim1_inst_MISO
		hps_io_hps_io_spim1_inst_SS0              : out   std_logic;                                        --                             .hps_io_spim1_inst_SS0
		hps_io_hps_io_uart0_inst_RX               : in    std_logic                     := '0';             --                             .hps_io_uart0_inst_RX
		hps_io_hps_io_uart0_inst_TX               : out   std_logic;                                        --                             .hps_io_uart0_inst_TX
		hps_io_hps_io_i2c0_inst_SDA               : inout std_logic                     := '0';             --                             .hps_io_i2c0_inst_SDA
		hps_io_hps_io_i2c0_inst_SCL               : inout std_logic                     := '0';             --                             .hps_io_i2c0_inst_SCL
		hps_io_hps_io_i2c1_inst_SDA               : inout std_logic                     := '0';             --                             .hps_io_i2c1_inst_SDA
		hps_io_hps_io_i2c1_inst_SCL               : inout std_logic                     := '0';             --                             .hps_io_i2c1_inst_SCL
		hps_io_hps_io_gpio_inst_GPIO09            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO09
		hps_io_hps_io_gpio_inst_GPIO35            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO35
		hps_io_hps_io_gpio_inst_GPIO37            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO37
		hps_io_hps_io_gpio_inst_GPIO40            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO40
		hps_io_hps_io_gpio_inst_GPIO41            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO41
		hps_io_hps_io_gpio_inst_GPIO44            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO44
		hps_io_hps_io_gpio_inst_GPIO48            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO48
		hps_io_hps_io_gpio_inst_GPIO53            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO53
		hps_io_hps_io_gpio_inst_GPIO54            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO54
		hps_io_hps_io_gpio_inst_GPIO61            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO61
		memory_mem_a                              : out   std_logic_vector(14 downto 0);                    --                       memory.mem_a
		memory_mem_ba                             : out   std_logic_vector(2 downto 0);                     --                             .mem_ba
		memory_mem_ck                             : out   std_logic;                                        --                             .mem_ck
		memory_mem_ck_n                           : out   std_logic;                                        --                             .mem_ck_n
		memory_mem_cke                            : out   std_logic;                                        --                             .mem_cke
		memory_mem_cs_n                           : out   std_logic;                                        --                             .mem_cs_n
		memory_mem_ras_n                          : out   std_logic;                                        --                             .mem_ras_n
		memory_mem_cas_n                          : out   std_logic;                                        --                             .mem_cas_n
		memory_mem_we_n                           : out   std_logic;                                        --                             .mem_we_n
		memory_mem_reset_n                        : out   std_logic;                                        --                             .mem_reset_n
		memory_mem_dq                             : inout std_logic_vector(31 downto 0) := (others => '0'); --                             .mem_dq
		memory_mem_dqs                            : inout std_logic_vector(3 downto 0)  := (others => '0'); --                             .mem_dqs
		memory_mem_dqs_n                          : inout std_logic_vector(3 downto 0)  := (others => '0'); --                             .mem_dqs_n
		memory_mem_odt                            : out   std_logic;                                        --                             .mem_odt
		memory_mem_dm                             : out   std_logic_vector(3 downto 0);                     --                             .mem_dm
		memory_oct_rzqin                          : in    std_logic                     := '0';             --                             .oct_rzqin
		sdram_addr                                : out   std_logic_vector(12 downto 0);                    --                        sdram.addr
		sdram_ba                                  : out   std_logic_vector(1 downto 0);                     --                             .ba
		sdram_cas_n                               : out   std_logic;                                        --                             .cas_n
		sdram_cke                                 : out   std_logic;                                        --                             .cke
		sdram_cs_n                                : out   std_logic;                                        --                             .cs_n
		sdram_dq                                  : inout std_logic_vector(15 downto 0) := (others => '0'); --                             .dq
		sdram_dqm                                 : out   std_logic_vector(1 downto 0);                     --                             .dqm
		sdram_ras_n                               : out   std_logic;                                        --                             .ras_n
		sdram_we_n                                : out   std_logic;                                        --                             .we_n
		system_pll_ref_clk_clk                    : in    std_logic                     := '0';             --           system_pll_ref_clk.clk
		system_pll_ref_reset_reset                : in    std_logic                     := '0'              --         system_pll_ref_reset.reset
	);
end entity dma_platform;

architecture rtl of dma_platform is
	component dma_platform_ARM_A9_HPS is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			f2h_stm_hwevents         : in    std_logic_vector(27 downto 0) := (others => 'X'); -- stm_hwevents
			mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                   : out   std_logic;                                        -- mem_ck
			mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
			mem_cke                  : out   std_logic;                                        -- mem_cke
			mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                : out   std_logic;                                        -- mem_cas_n
			mem_we_n                 : out   std_logic;                                        -- mem_we_n
			mem_reset_n              : out   std_logic;                                        -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                        -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_qspi_inst_IO0     : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO0
			hps_io_qspi_inst_IO1     : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO1
			hps_io_qspi_inst_IO2     : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO2
			hps_io_qspi_inst_IO3     : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO3
			hps_io_qspi_inst_SS0     : out   std_logic;                                        -- hps_io_qspi_inst_SS0
			hps_io_qspi_inst_CLK     : out   std_logic;                                        -- hps_io_qspi_inst_CLK
			hps_io_sdio_inst_CMD     : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                        -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim0_inst_CLK    : out   std_logic;                                        -- hps_io_spim0_inst_CLK
			hps_io_spim0_inst_MOSI   : out   std_logic;                                        -- hps_io_spim0_inst_MOSI
			hps_io_spim0_inst_MISO   : in    std_logic                     := 'X';             -- hps_io_spim0_inst_MISO
			hps_io_spim0_inst_SS0    : out   std_logic;                                        -- hps_io_spim0_inst_SS0
			hps_io_spim1_inst_CLK    : out   std_logic;                                        -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   : out   std_logic;                                        -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   : in    std_logic                     := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    : out   std_logic;                                        -- hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO37  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO37
			hps_io_gpio_inst_GPIO40  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO41  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO41
			hps_io_gpio_inst_GPIO44  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO44
			hps_io_gpio_inst_GPIO48  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO61
			h2f_rst_n                : out   std_logic;                                        -- reset_n
			h2f_axi_clk              : in    std_logic                     := 'X';             -- clk
			h2f_AWID                 : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_AWADDR               : out   std_logic_vector(29 downto 0);                    -- awaddr
			h2f_AWLEN                : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_AWSIZE               : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_AWBURST              : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_AWLOCK               : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_AWCACHE              : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_AWPROT               : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_AWVALID              : out   std_logic;                                        -- awvalid
			h2f_AWREADY              : in    std_logic                     := 'X';             -- awready
			h2f_WID                  : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_WDATA                : out   std_logic_vector(63 downto 0);                    -- wdata
			h2f_WSTRB                : out   std_logic_vector(7 downto 0);                     -- wstrb
			h2f_WLAST                : out   std_logic;                                        -- wlast
			h2f_WVALID               : out   std_logic;                                        -- wvalid
			h2f_WREADY               : in    std_logic                     := 'X';             -- wready
			h2f_BID                  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_BRESP                : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_BVALID               : in    std_logic                     := 'X';             -- bvalid
			h2f_BREADY               : out   std_logic;                                        -- bready
			h2f_ARID                 : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_ARADDR               : out   std_logic_vector(29 downto 0);                    -- araddr
			h2f_ARLEN                : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_ARSIZE               : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_ARBURST              : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_ARLOCK               : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_ARCACHE              : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_ARPROT               : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_ARVALID              : out   std_logic;                                        -- arvalid
			h2f_ARREADY              : in    std_logic                     := 'X';             -- arready
			h2f_RID                  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_RDATA                : in    std_logic_vector(63 downto 0) := (others => 'X'); -- rdata
			h2f_RRESP                : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_RLAST                : in    std_logic                     := 'X';             -- rlast
			h2f_RVALID               : in    std_logic                     := 'X';             -- rvalid
			h2f_RREADY               : out   std_logic;                                        -- rready
			f2h_axi_clk              : in    std_logic                     := 'X';             -- clk
			f2h_AWID                 : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- awid
			f2h_AWADDR               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			f2h_AWLEN                : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			f2h_AWSIZE               : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			f2h_AWBURST              : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			f2h_AWLOCK               : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			f2h_AWCACHE              : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			f2h_AWPROT               : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			f2h_AWVALID              : in    std_logic                     := 'X';             -- awvalid
			f2h_AWREADY              : out   std_logic;                                        -- awready
			f2h_AWUSER               : in    std_logic_vector(4 downto 0)  := (others => 'X'); -- awuser
			f2h_WID                  : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- wid
			f2h_WDATA                : in    std_logic_vector(63 downto 0) := (others => 'X'); -- wdata
			f2h_WSTRB                : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- wstrb
			f2h_WLAST                : in    std_logic                     := 'X';             -- wlast
			f2h_WVALID               : in    std_logic                     := 'X';             -- wvalid
			f2h_WREADY               : out   std_logic;                                        -- wready
			f2h_BID                  : out   std_logic_vector(7 downto 0);                     -- bid
			f2h_BRESP                : out   std_logic_vector(1 downto 0);                     -- bresp
			f2h_BVALID               : out   std_logic;                                        -- bvalid
			f2h_BREADY               : in    std_logic                     := 'X';             -- bready
			f2h_ARID                 : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- arid
			f2h_ARADDR               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			f2h_ARLEN                : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			f2h_ARSIZE               : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			f2h_ARBURST              : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			f2h_ARLOCK               : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			f2h_ARCACHE              : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			f2h_ARPROT               : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			f2h_ARVALID              : in    std_logic                     := 'X';             -- arvalid
			f2h_ARREADY              : out   std_logic;                                        -- arready
			f2h_ARUSER               : in    std_logic_vector(4 downto 0)  := (others => 'X'); -- aruser
			f2h_RID                  : out   std_logic_vector(7 downto 0);                     -- rid
			f2h_RDATA                : out   std_logic_vector(63 downto 0);                    -- rdata
			f2h_RRESP                : out   std_logic_vector(1 downto 0);                     -- rresp
			f2h_RLAST                : out   std_logic;                                        -- rlast
			f2h_RVALID               : out   std_logic;                                        -- rvalid
			f2h_RREADY               : in    std_logic                     := 'X';             -- rready
			h2f_lw_axi_clk           : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY           : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                        -- wlast
			h2f_lw_WVALID            : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY            : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                        -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY           : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic;                                        -- rready
			f2h_irq_p0               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			f2h_irq_p1               : in    std_logic_vector(31 downto 0) := (others => 'X')  -- irq
		);
	end component dma_platform_ARM_A9_HPS;

	component anomaly_detection is
		generic (
			IM_SIZE     : integer := 500;
			ADDR_SIZE   : integer := 16;
			WORD_SIZE   : integer := 16;
			COUNT_WIDTH : integer := 9
		);
		port (
			clk             : in  std_logic                     := 'X';             -- clk
			rst             : in  std_logic                     := 'X';             -- reset
			data_out        : out std_logic_vector(15 downto 0);                    -- data
			endpacket_out   : out std_logic;                                        -- endofpacket
			ready_in        : in  std_logic                     := 'X';             -- ready
			startpacket_out : out std_logic;                                        -- startofpacket
			valid_out       : out std_logic;                                        -- valid
			data_in         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			endpacket_in    : in  std_logic                     := 'X';             -- endofpacket
			ready_out       : out std_logic;                                        -- ready
			startpacket_in  : in  std_logic                     := 'X';             -- startofpacket
			valid_in        : in  std_logic                     := 'X'              -- valid
		);
	end component anomaly_detection;

	component dma_platform_Change_Detection_Mem_to_Stream_DMA is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_data          : out std_logic_vector(15 downto 0);                    -- data
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic                                         -- valid
		);
	end component dma_platform_Change_Detection_Mem_to_Stream_DMA;

	component altera_up_avalon_video_dma_ctrl_addr_trans is
		generic (
			ADDRESS_TRANSLATION_MASK : std_logic_vector(31 downto 0) := "11000000000000000000000000000000"
		);
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			slave_address      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read         : in  std_logic                     := 'X';             -- read
			slave_write        : in  std_logic                     := 'X';             -- write
			slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			slave_waitrequest  : out std_logic;                                        -- waitrequest
			master_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			master_address     : out std_logic_vector(1 downto 0);                     -- address
			master_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			master_read        : out std_logic;                                        -- read
			master_write       : out std_logic;                                        -- write
			master_writedata   : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component altera_up_avalon_video_dma_ctrl_addr_trans;

	component dma_platform_Change_Detection_Stream_to_Mem_DMA is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			stream_data          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			stream_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			stream_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			stream_valid         : in  std_logic                     := 'X';             -- valid
			stream_ready         : out std_logic;                                        -- ready
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(15 downto 0)                     -- writedata
		);
	end component dma_platform_Change_Detection_Stream_to_Mem_DMA;

	component dma_platform_SDRAM is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component dma_platform_SDRAM;

	component dma_platform_System_PLL is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component dma_platform_System_PLL;

	component dma_platform_mm_interconnect_0 is
		port (
			ARM_A9_HPS_h2f_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			ARM_A9_HPS_h2f_axi_master_awaddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- awaddr
			ARM_A9_HPS_h2f_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			ARM_A9_HPS_h2f_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			ARM_A9_HPS_h2f_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			ARM_A9_HPS_h2f_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			ARM_A9_HPS_h2f_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			ARM_A9_HPS_h2f_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			ARM_A9_HPS_h2f_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			ARM_A9_HPS_h2f_axi_master_awready                                     : out std_logic;                                        -- awready
			ARM_A9_HPS_h2f_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			ARM_A9_HPS_h2f_axi_master_wdata                                       : in  std_logic_vector(63 downto 0) := (others => 'X'); -- wdata
			ARM_A9_HPS_h2f_axi_master_wstrb                                       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wstrb
			ARM_A9_HPS_h2f_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			ARM_A9_HPS_h2f_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			ARM_A9_HPS_h2f_axi_master_wready                                      : out std_logic;                                        -- wready
			ARM_A9_HPS_h2f_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			ARM_A9_HPS_h2f_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			ARM_A9_HPS_h2f_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			ARM_A9_HPS_h2f_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			ARM_A9_HPS_h2f_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			ARM_A9_HPS_h2f_axi_master_araddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- araddr
			ARM_A9_HPS_h2f_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			ARM_A9_HPS_h2f_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			ARM_A9_HPS_h2f_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			ARM_A9_HPS_h2f_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			ARM_A9_HPS_h2f_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			ARM_A9_HPS_h2f_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			ARM_A9_HPS_h2f_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			ARM_A9_HPS_h2f_axi_master_arready                                     : out std_logic;                                        -- arready
			ARM_A9_HPS_h2f_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			ARM_A9_HPS_h2f_axi_master_rdata                                       : out std_logic_vector(63 downto 0);                    -- rdata
			ARM_A9_HPS_h2f_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			ARM_A9_HPS_h2f_axi_master_rlast                                       : out std_logic;                                        -- rlast
			ARM_A9_HPS_h2f_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			ARM_A9_HPS_h2f_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			System_PLL_sys_clk_clk                                                : in  std_logic                     := 'X';             -- clk
			ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Change_Detection_Mem_to_Stream_DMA_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_address          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_waitrequest      : out std_logic;                                        -- waitrequest
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_read             : in  std_logic                     := 'X';             -- read
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_readdata         : out std_logic_vector(15 downto 0);                    -- readdata
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_readdatavalid    : out std_logic;                                        -- readdatavalid
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_lock             : in  std_logic                     := 'X';             -- lock
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_master_address          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_master_waitrequest      : out std_logic;                                        -- waitrequest
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_master_write            : in  std_logic                     := 'X';             -- write
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_master_writedata        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			SDRAM_s1_address                                                      : out std_logic_vector(24 downto 0);                    -- address
			SDRAM_s1_write                                                        : out std_logic;                                        -- write
			SDRAM_s1_read                                                         : out std_logic;                                        -- read
			SDRAM_s1_readdata                                                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SDRAM_s1_writedata                                                    : out std_logic_vector(15 downto 0);                    -- writedata
			SDRAM_s1_byteenable                                                   : out std_logic_vector(1 downto 0);                     -- byteenable
			SDRAM_s1_readdatavalid                                                : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_s1_waitrequest                                                  : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_s1_chipselect                                                   : out std_logic                                         -- chipselect
		);
	end component dma_platform_mm_interconnect_0;

	component dma_platform_mm_interconnect_1 is
		port (
			ARM_A9_HPS_h2f_lw_axi_master_awid                                           : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			ARM_A9_HPS_h2f_lw_axi_master_awaddr                                         : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			ARM_A9_HPS_h2f_lw_axi_master_awlen                                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			ARM_A9_HPS_h2f_lw_axi_master_awsize                                         : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			ARM_A9_HPS_h2f_lw_axi_master_awburst                                        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			ARM_A9_HPS_h2f_lw_axi_master_awlock                                         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			ARM_A9_HPS_h2f_lw_axi_master_awcache                                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			ARM_A9_HPS_h2f_lw_axi_master_awprot                                         : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			ARM_A9_HPS_h2f_lw_axi_master_awvalid                                        : in  std_logic                     := 'X';             -- awvalid
			ARM_A9_HPS_h2f_lw_axi_master_awready                                        : out std_logic;                                        -- awready
			ARM_A9_HPS_h2f_lw_axi_master_wid                                            : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			ARM_A9_HPS_h2f_lw_axi_master_wdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			ARM_A9_HPS_h2f_lw_axi_master_wstrb                                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			ARM_A9_HPS_h2f_lw_axi_master_wlast                                          : in  std_logic                     := 'X';             -- wlast
			ARM_A9_HPS_h2f_lw_axi_master_wvalid                                         : in  std_logic                     := 'X';             -- wvalid
			ARM_A9_HPS_h2f_lw_axi_master_wready                                         : out std_logic;                                        -- wready
			ARM_A9_HPS_h2f_lw_axi_master_bid                                            : out std_logic_vector(11 downto 0);                    -- bid
			ARM_A9_HPS_h2f_lw_axi_master_bresp                                          : out std_logic_vector(1 downto 0);                     -- bresp
			ARM_A9_HPS_h2f_lw_axi_master_bvalid                                         : out std_logic;                                        -- bvalid
			ARM_A9_HPS_h2f_lw_axi_master_bready                                         : in  std_logic                     := 'X';             -- bready
			ARM_A9_HPS_h2f_lw_axi_master_arid                                           : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			ARM_A9_HPS_h2f_lw_axi_master_araddr                                         : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			ARM_A9_HPS_h2f_lw_axi_master_arlen                                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			ARM_A9_HPS_h2f_lw_axi_master_arsize                                         : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			ARM_A9_HPS_h2f_lw_axi_master_arburst                                        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			ARM_A9_HPS_h2f_lw_axi_master_arlock                                         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			ARM_A9_HPS_h2f_lw_axi_master_arcache                                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			ARM_A9_HPS_h2f_lw_axi_master_arprot                                         : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			ARM_A9_HPS_h2f_lw_axi_master_arvalid                                        : in  std_logic                     := 'X';             -- arvalid
			ARM_A9_HPS_h2f_lw_axi_master_arready                                        : out std_logic;                                        -- arready
			ARM_A9_HPS_h2f_lw_axi_master_rid                                            : out std_logic_vector(11 downto 0);                    -- rid
			ARM_A9_HPS_h2f_lw_axi_master_rdata                                          : out std_logic_vector(31 downto 0);                    -- rdata
			ARM_A9_HPS_h2f_lw_axi_master_rresp                                          : out std_logic_vector(1 downto 0);                     -- rresp
			ARM_A9_HPS_h2f_lw_axi_master_rlast                                          : out std_logic;                                        -- rlast
			ARM_A9_HPS_h2f_lw_axi_master_rvalid                                         : out std_logic;                                        -- rvalid
			ARM_A9_HPS_h2f_lw_axi_master_rready                                         : in  std_logic                     := 'X';             -- rready
			System_PLL_sys_clk_clk                                                      : in  std_logic                     := 'X';             -- clk
			ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset    : in  std_logic                     := 'X';             -- reset
			Change_Detection_Mem_to_Stream_Translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Change_Detection_Mem_to_Stream_Translator_slave_address                     : out std_logic_vector(1 downto 0);                     -- address
			Change_Detection_Mem_to_Stream_Translator_slave_write                       : out std_logic;                                        -- write
			Change_Detection_Mem_to_Stream_Translator_slave_read                        : out std_logic;                                        -- read
			Change_Detection_Mem_to_Stream_Translator_slave_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Change_Detection_Mem_to_Stream_Translator_slave_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			Change_Detection_Mem_to_Stream_Translator_slave_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			Change_Detection_Mem_to_Stream_Translator_slave_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			Change_Detection_Stream_to_Mem_Translator_slave_address                     : out std_logic_vector(1 downto 0);                     -- address
			Change_Detection_Stream_to_Mem_Translator_slave_write                       : out std_logic;                                        -- write
			Change_Detection_Stream_to_Mem_Translator_slave_read                        : out std_logic;                                        -- read
			Change_Detection_Stream_to_Mem_Translator_slave_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Change_Detection_Stream_to_Mem_Translator_slave_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			Change_Detection_Stream_to_Mem_Translator_slave_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			Change_Detection_Stream_to_Mem_Translator_slave_waitrequest                 : in  std_logic                     := 'X'              -- waitrequest
		);
	end component dma_platform_mm_interconnect_1;

	component dma_platform_mm_interconnect_2 is
		port (
			System_PLL_sys_clk_clk                                                      : in  std_logic                     := 'X';             -- clk
			Change_Detection_Mem_to_Stream_Translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Change_Detection_Mem_to_Stream_Translator_master_address                    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			Change_Detection_Mem_to_Stream_Translator_master_waitrequest                : out std_logic;                                        -- waitrequest
			Change_Detection_Mem_to_Stream_Translator_master_byteenable                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Change_Detection_Mem_to_Stream_Translator_master_read                       : in  std_logic                     := 'X';             -- read
			Change_Detection_Mem_to_Stream_Translator_master_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			Change_Detection_Mem_to_Stream_Translator_master_write                      : in  std_logic                     := 'X';             -- write
			Change_Detection_Mem_to_Stream_Translator_master_writedata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_address         : out std_logic_vector(1 downto 0);                     -- address
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_write           : out std_logic;                                        -- write
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_read            : out std_logic;                                        -- read
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_writedata       : out std_logic_vector(31 downto 0);                    -- writedata
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_byteenable      : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component dma_platform_mm_interconnect_2;

	component dma_platform_mm_interconnect_3 is
		port (
			System_PLL_sys_clk_clk                                                      : in  std_logic                     := 'X';             -- clk
			Change_Detection_Stream_to_Mem_Translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Change_Detection_Stream_to_Mem_Translator_master_address                    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			Change_Detection_Stream_to_Mem_Translator_master_waitrequest                : out std_logic;                                        -- waitrequest
			Change_Detection_Stream_to_Mem_Translator_master_byteenable                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Change_Detection_Stream_to_Mem_Translator_master_read                       : in  std_logic                     := 'X';             -- read
			Change_Detection_Stream_to_Mem_Translator_master_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			Change_Detection_Stream_to_Mem_Translator_master_write                      : in  std_logic                     := 'X';             -- write
			Change_Detection_Stream_to_Mem_Translator_master_writedata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_address         : out std_logic_vector(1 downto 0);                     -- address
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_write           : out std_logic;                                        -- write
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_read            : out std_logic;                                        -- read
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_writedata       : out std_logic_vector(31 downto 0);                    -- writedata
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_byteenable      : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component dma_platform_mm_interconnect_3;

	component dma_platform_irq_mapper is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component dma_platform_irq_mapper;

	component dma_platform_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component dma_platform_rst_controller;

	component dma_platform_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component dma_platform_rst_controller_001;

	signal change_detection_mem_to_stream_dma_avalon_pixel_source_valid                             : std_logic;                     -- Change_Detection_Mem_to_Stream_DMA:stream_valid -> Anomaly_Detection_Module:valid_in
	signal change_detection_mem_to_stream_dma_avalon_pixel_source_data                              : std_logic_vector(15 downto 0); -- Change_Detection_Mem_to_Stream_DMA:stream_data -> Anomaly_Detection_Module:data_in
	signal change_detection_mem_to_stream_dma_avalon_pixel_source_ready                             : std_logic;                     -- Anomaly_Detection_Module:ready_out -> Change_Detection_Mem_to_Stream_DMA:stream_ready
	signal change_detection_mem_to_stream_dma_avalon_pixel_source_startofpacket                     : std_logic;                     -- Change_Detection_Mem_to_Stream_DMA:stream_startofpacket -> Anomaly_Detection_Module:startpacket_in
	signal change_detection_mem_to_stream_dma_avalon_pixel_source_endofpacket                       : std_logic;                     -- Change_Detection_Mem_to_Stream_DMA:stream_endofpacket -> Anomaly_Detection_Module:endpacket_in
	signal anomaly_detection_module_avalon_streaming_source_valid                                   : std_logic;                     -- Anomaly_Detection_Module:valid_out -> Change_Detection_Stream_to_Mem_DMA:stream_valid
	signal anomaly_detection_module_avalon_streaming_source_data                                    : std_logic_vector(15 downto 0); -- Anomaly_Detection_Module:data_out -> Change_Detection_Stream_to_Mem_DMA:stream_data
	signal anomaly_detection_module_avalon_streaming_source_ready                                   : std_logic;                     -- Change_Detection_Stream_to_Mem_DMA:stream_ready -> Anomaly_Detection_Module:ready_in
	signal anomaly_detection_module_avalon_streaming_source_startofpacket                           : std_logic;                     -- Anomaly_Detection_Module:startpacket_out -> Change_Detection_Stream_to_Mem_DMA:stream_startofpacket
	signal anomaly_detection_module_avalon_streaming_source_endofpacket                             : std_logic;                     -- Anomaly_Detection_Module:endpacket_out -> Change_Detection_Stream_to_Mem_DMA:stream_endofpacket
	signal system_pll_sys_clk_clk                                                                   : std_logic;                     -- System_PLL:sys_clk_clk -> [ARM_A9_HPS:f2h_axi_clk, ARM_A9_HPS:h2f_axi_clk, ARM_A9_HPS:h2f_lw_axi_clk, Anomaly_Detection_Module:clk, Change_Detection_Mem_to_Stream_DMA:clk, Change_Detection_Mem_to_Stream_Translator:clk, Change_Detection_Stream_to_Mem_DMA:clk, Change_Detection_Stream_to_Mem_Translator:clk, SDRAM:clk, mm_interconnect_0:System_PLL_sys_clk_clk, mm_interconnect_1:System_PLL_sys_clk_clk, mm_interconnect_2:System_PLL_sys_clk_clk, mm_interconnect_3:System_PLL_sys_clk_clk, rst_controller:clk, rst_controller_001:clk]
	signal change_detection_mem_to_stream_dma_avalon_dma_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_waitrequest -> Change_Detection_Mem_to_Stream_DMA:master_waitrequest
	signal change_detection_mem_to_stream_dma_avalon_dma_master_readdata                            : std_logic_vector(15 downto 0); -- mm_interconnect_0:Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_readdata -> Change_Detection_Mem_to_Stream_DMA:master_readdata
	signal change_detection_mem_to_stream_dma_avalon_dma_master_address                             : std_logic_vector(31 downto 0); -- Change_Detection_Mem_to_Stream_DMA:master_address -> mm_interconnect_0:Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_address
	signal change_detection_mem_to_stream_dma_avalon_dma_master_read                                : std_logic;                     -- Change_Detection_Mem_to_Stream_DMA:master_read -> mm_interconnect_0:Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_read
	signal change_detection_mem_to_stream_dma_avalon_dma_master_readdatavalid                       : std_logic;                     -- mm_interconnect_0:Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_readdatavalid -> Change_Detection_Mem_to_Stream_DMA:master_readdatavalid
	signal change_detection_mem_to_stream_dma_avalon_dma_master_lock                                : std_logic;                     -- Change_Detection_Mem_to_Stream_DMA:master_arbiterlock -> mm_interconnect_0:Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_lock
	signal change_detection_stream_to_mem_dma_avalon_dma_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:Change_Detection_Stream_to_Mem_DMA_avalon_dma_master_waitrequest -> Change_Detection_Stream_to_Mem_DMA:master_waitrequest
	signal change_detection_stream_to_mem_dma_avalon_dma_master_address                             : std_logic_vector(31 downto 0); -- Change_Detection_Stream_to_Mem_DMA:master_address -> mm_interconnect_0:Change_Detection_Stream_to_Mem_DMA_avalon_dma_master_address
	signal change_detection_stream_to_mem_dma_avalon_dma_master_write                               : std_logic;                     -- Change_Detection_Stream_to_Mem_DMA:master_write -> mm_interconnect_0:Change_Detection_Stream_to_Mem_DMA_avalon_dma_master_write
	signal change_detection_stream_to_mem_dma_avalon_dma_master_writedata                           : std_logic_vector(15 downto 0); -- Change_Detection_Stream_to_Mem_DMA:master_writedata -> mm_interconnect_0:Change_Detection_Stream_to_Mem_DMA_avalon_dma_master_writedata
	signal arm_a9_hps_h2f_axi_master_awburst                                                        : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_AWBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awburst
	signal arm_a9_hps_h2f_axi_master_arlen                                                          : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_ARLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlen
	signal arm_a9_hps_h2f_axi_master_wstrb                                                          : std_logic_vector(7 downto 0);  -- ARM_A9_HPS:h2f_WSTRB -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wstrb
	signal arm_a9_hps_h2f_axi_master_wready                                                         : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wready -> ARM_A9_HPS:h2f_WREADY
	signal arm_a9_hps_h2f_axi_master_rid                                                            : std_logic_vector(11 downto 0); -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rid -> ARM_A9_HPS:h2f_RID
	signal arm_a9_hps_h2f_axi_master_rready                                                         : std_logic;                     -- ARM_A9_HPS:h2f_RREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rready
	signal arm_a9_hps_h2f_axi_master_awlen                                                          : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_AWLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlen
	signal arm_a9_hps_h2f_axi_master_wid                                                            : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_WID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wid
	signal arm_a9_hps_h2f_axi_master_arcache                                                        : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_ARCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arcache
	signal arm_a9_hps_h2f_axi_master_wvalid                                                         : std_logic;                     -- ARM_A9_HPS:h2f_WVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wvalid
	signal arm_a9_hps_h2f_axi_master_araddr                                                         : std_logic_vector(29 downto 0); -- ARM_A9_HPS:h2f_ARADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_araddr
	signal arm_a9_hps_h2f_axi_master_arprot                                                         : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_ARPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arprot
	signal arm_a9_hps_h2f_axi_master_awprot                                                         : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_AWPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awprot
	signal arm_a9_hps_h2f_axi_master_wdata                                                          : std_logic_vector(63 downto 0); -- ARM_A9_HPS:h2f_WDATA -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wdata
	signal arm_a9_hps_h2f_axi_master_arvalid                                                        : std_logic;                     -- ARM_A9_HPS:h2f_ARVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arvalid
	signal arm_a9_hps_h2f_axi_master_awcache                                                        : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_AWCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awcache
	signal arm_a9_hps_h2f_axi_master_arid                                                           : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_ARID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arid
	signal arm_a9_hps_h2f_axi_master_arlock                                                         : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_ARLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlock
	signal arm_a9_hps_h2f_axi_master_awlock                                                         : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_AWLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlock
	signal arm_a9_hps_h2f_axi_master_awaddr                                                         : std_logic_vector(29 downto 0); -- ARM_A9_HPS:h2f_AWADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awaddr
	signal arm_a9_hps_h2f_axi_master_bresp                                                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bresp -> ARM_A9_HPS:h2f_BRESP
	signal arm_a9_hps_h2f_axi_master_arready                                                        : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arready -> ARM_A9_HPS:h2f_ARREADY
	signal arm_a9_hps_h2f_axi_master_rdata                                                          : std_logic_vector(63 downto 0); -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rdata -> ARM_A9_HPS:h2f_RDATA
	signal arm_a9_hps_h2f_axi_master_awready                                                        : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awready -> ARM_A9_HPS:h2f_AWREADY
	signal arm_a9_hps_h2f_axi_master_arburst                                                        : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_ARBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arburst
	signal arm_a9_hps_h2f_axi_master_arsize                                                         : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_ARSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arsize
	signal arm_a9_hps_h2f_axi_master_bready                                                         : std_logic;                     -- ARM_A9_HPS:h2f_BREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bready
	signal arm_a9_hps_h2f_axi_master_rlast                                                          : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rlast -> ARM_A9_HPS:h2f_RLAST
	signal arm_a9_hps_h2f_axi_master_wlast                                                          : std_logic;                     -- ARM_A9_HPS:h2f_WLAST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wlast
	signal arm_a9_hps_h2f_axi_master_rresp                                                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rresp -> ARM_A9_HPS:h2f_RRESP
	signal arm_a9_hps_h2f_axi_master_awid                                                           : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_AWID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awid
	signal arm_a9_hps_h2f_axi_master_bid                                                            : std_logic_vector(11 downto 0); -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bid -> ARM_A9_HPS:h2f_BID
	signal arm_a9_hps_h2f_axi_master_bvalid                                                         : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bvalid -> ARM_A9_HPS:h2f_BVALID
	signal arm_a9_hps_h2f_axi_master_awsize                                                         : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_AWSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awsize
	signal arm_a9_hps_h2f_axi_master_awvalid                                                        : std_logic;                     -- ARM_A9_HPS:h2f_AWVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awvalid
	signal arm_a9_hps_h2f_axi_master_rvalid                                                         : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rvalid -> ARM_A9_HPS:h2f_RVALID
	signal mm_interconnect_0_sdram_s1_chipselect                                                    : std_logic;                     -- mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                                                      : std_logic_vector(15 downto 0); -- SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                                                   : std_logic;                     -- SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                                       : std_logic_vector(24 downto 0); -- mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	signal mm_interconnect_0_sdram_s1_read                                                          : std_logic;                     -- mm_interconnect_0:SDRAM_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SDRAM_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                                                 : std_logic;                     -- SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                                         : std_logic;                     -- mm_interconnect_0:SDRAM_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                                                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	signal arm_a9_hps_h2f_lw_axi_master_awburst                                                     : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_lw_AWBURST -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awburst
	signal arm_a9_hps_h2f_lw_axi_master_arlen                                                       : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_ARLEN -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arlen
	signal arm_a9_hps_h2f_lw_axi_master_wstrb                                                       : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_WSTRB -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wstrb
	signal arm_a9_hps_h2f_lw_axi_master_wready                                                      : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wready -> ARM_A9_HPS:h2f_lw_WREADY
	signal arm_a9_hps_h2f_lw_axi_master_rid                                                         : std_logic_vector(11 downto 0); -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rid -> ARM_A9_HPS:h2f_lw_RID
	signal arm_a9_hps_h2f_lw_axi_master_rready                                                      : std_logic;                     -- ARM_A9_HPS:h2f_lw_RREADY -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rready
	signal arm_a9_hps_h2f_lw_axi_master_awlen                                                       : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_AWLEN -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awlen
	signal arm_a9_hps_h2f_lw_axi_master_wid                                                         : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_lw_WID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wid
	signal arm_a9_hps_h2f_lw_axi_master_arcache                                                     : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_ARCACHE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arcache
	signal arm_a9_hps_h2f_lw_axi_master_wvalid                                                      : std_logic;                     -- ARM_A9_HPS:h2f_lw_WVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wvalid
	signal arm_a9_hps_h2f_lw_axi_master_araddr                                                      : std_logic_vector(20 downto 0); -- ARM_A9_HPS:h2f_lw_ARADDR -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_araddr
	signal arm_a9_hps_h2f_lw_axi_master_arprot                                                      : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_lw_ARPROT -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arprot
	signal arm_a9_hps_h2f_lw_axi_master_awprot                                                      : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_lw_AWPROT -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awprot
	signal arm_a9_hps_h2f_lw_axi_master_wdata                                                       : std_logic_vector(31 downto 0); -- ARM_A9_HPS:h2f_lw_WDATA -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wdata
	signal arm_a9_hps_h2f_lw_axi_master_arvalid                                                     : std_logic;                     -- ARM_A9_HPS:h2f_lw_ARVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arvalid
	signal arm_a9_hps_h2f_lw_axi_master_awcache                                                     : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_AWCACHE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awcache
	signal arm_a9_hps_h2f_lw_axi_master_arid                                                        : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_lw_ARID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arid
	signal arm_a9_hps_h2f_lw_axi_master_arlock                                                      : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_lw_ARLOCK -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arlock
	signal arm_a9_hps_h2f_lw_axi_master_awlock                                                      : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_lw_AWLOCK -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awlock
	signal arm_a9_hps_h2f_lw_axi_master_awaddr                                                      : std_logic_vector(20 downto 0); -- ARM_A9_HPS:h2f_lw_AWADDR -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awaddr
	signal arm_a9_hps_h2f_lw_axi_master_bresp                                                       : std_logic_vector(1 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bresp -> ARM_A9_HPS:h2f_lw_BRESP
	signal arm_a9_hps_h2f_lw_axi_master_arready                                                     : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arready -> ARM_A9_HPS:h2f_lw_ARREADY
	signal arm_a9_hps_h2f_lw_axi_master_rdata                                                       : std_logic_vector(31 downto 0); -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rdata -> ARM_A9_HPS:h2f_lw_RDATA
	signal arm_a9_hps_h2f_lw_axi_master_awready                                                     : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awready -> ARM_A9_HPS:h2f_lw_AWREADY
	signal arm_a9_hps_h2f_lw_axi_master_arburst                                                     : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_lw_ARBURST -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arburst
	signal arm_a9_hps_h2f_lw_axi_master_arsize                                                      : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_lw_ARSIZE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arsize
	signal arm_a9_hps_h2f_lw_axi_master_bready                                                      : std_logic;                     -- ARM_A9_HPS:h2f_lw_BREADY -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bready
	signal arm_a9_hps_h2f_lw_axi_master_rlast                                                       : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rlast -> ARM_A9_HPS:h2f_lw_RLAST
	signal arm_a9_hps_h2f_lw_axi_master_wlast                                                       : std_logic;                     -- ARM_A9_HPS:h2f_lw_WLAST -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wlast
	signal arm_a9_hps_h2f_lw_axi_master_rresp                                                       : std_logic_vector(1 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rresp -> ARM_A9_HPS:h2f_lw_RRESP
	signal arm_a9_hps_h2f_lw_axi_master_awid                                                        : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_lw_AWID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awid
	signal arm_a9_hps_h2f_lw_axi_master_bid                                                         : std_logic_vector(11 downto 0); -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bid -> ARM_A9_HPS:h2f_lw_BID
	signal arm_a9_hps_h2f_lw_axi_master_bvalid                                                      : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bvalid -> ARM_A9_HPS:h2f_lw_BVALID
	signal arm_a9_hps_h2f_lw_axi_master_awsize                                                      : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_lw_AWSIZE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awsize
	signal arm_a9_hps_h2f_lw_axi_master_awvalid                                                     : std_logic;                     -- ARM_A9_HPS:h2f_lw_AWVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awvalid
	signal arm_a9_hps_h2f_lw_axi_master_rvalid                                                      : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rvalid -> ARM_A9_HPS:h2f_lw_RVALID
	signal mm_interconnect_1_change_detection_mem_to_stream_translator_slave_readdata               : std_logic_vector(31 downto 0); -- Change_Detection_Mem_to_Stream_Translator:slave_readdata -> mm_interconnect_1:Change_Detection_Mem_to_Stream_Translator_slave_readdata
	signal mm_interconnect_1_change_detection_mem_to_stream_translator_slave_waitrequest            : std_logic;                     -- Change_Detection_Mem_to_Stream_Translator:slave_waitrequest -> mm_interconnect_1:Change_Detection_Mem_to_Stream_Translator_slave_waitrequest
	signal mm_interconnect_1_change_detection_mem_to_stream_translator_slave_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_1:Change_Detection_Mem_to_Stream_Translator_slave_address -> Change_Detection_Mem_to_Stream_Translator:slave_address
	signal mm_interconnect_1_change_detection_mem_to_stream_translator_slave_read                   : std_logic;                     -- mm_interconnect_1:Change_Detection_Mem_to_Stream_Translator_slave_read -> Change_Detection_Mem_to_Stream_Translator:slave_read
	signal mm_interconnect_1_change_detection_mem_to_stream_translator_slave_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_1:Change_Detection_Mem_to_Stream_Translator_slave_byteenable -> Change_Detection_Mem_to_Stream_Translator:slave_byteenable
	signal mm_interconnect_1_change_detection_mem_to_stream_translator_slave_write                  : std_logic;                     -- mm_interconnect_1:Change_Detection_Mem_to_Stream_Translator_slave_write -> Change_Detection_Mem_to_Stream_Translator:slave_write
	signal mm_interconnect_1_change_detection_mem_to_stream_translator_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_1:Change_Detection_Mem_to_Stream_Translator_slave_writedata -> Change_Detection_Mem_to_Stream_Translator:slave_writedata
	signal mm_interconnect_1_change_detection_stream_to_mem_translator_slave_readdata               : std_logic_vector(31 downto 0); -- Change_Detection_Stream_to_Mem_Translator:slave_readdata -> mm_interconnect_1:Change_Detection_Stream_to_Mem_Translator_slave_readdata
	signal mm_interconnect_1_change_detection_stream_to_mem_translator_slave_waitrequest            : std_logic;                     -- Change_Detection_Stream_to_Mem_Translator:slave_waitrequest -> mm_interconnect_1:Change_Detection_Stream_to_Mem_Translator_slave_waitrequest
	signal mm_interconnect_1_change_detection_stream_to_mem_translator_slave_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_1:Change_Detection_Stream_to_Mem_Translator_slave_address -> Change_Detection_Stream_to_Mem_Translator:slave_address
	signal mm_interconnect_1_change_detection_stream_to_mem_translator_slave_read                   : std_logic;                     -- mm_interconnect_1:Change_Detection_Stream_to_Mem_Translator_slave_read -> Change_Detection_Stream_to_Mem_Translator:slave_read
	signal mm_interconnect_1_change_detection_stream_to_mem_translator_slave_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_1:Change_Detection_Stream_to_Mem_Translator_slave_byteenable -> Change_Detection_Stream_to_Mem_Translator:slave_byteenable
	signal mm_interconnect_1_change_detection_stream_to_mem_translator_slave_write                  : std_logic;                     -- mm_interconnect_1:Change_Detection_Stream_to_Mem_Translator_slave_write -> Change_Detection_Stream_to_Mem_Translator:slave_write
	signal mm_interconnect_1_change_detection_stream_to_mem_translator_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_1:Change_Detection_Stream_to_Mem_Translator_slave_writedata -> Change_Detection_Stream_to_Mem_Translator:slave_writedata
	signal change_detection_mem_to_stream_translator_master_readdata                                : std_logic_vector(31 downto 0); -- mm_interconnect_2:Change_Detection_Mem_to_Stream_Translator_master_readdata -> Change_Detection_Mem_to_Stream_Translator:master_readdata
	signal change_detection_mem_to_stream_translator_master_waitrequest                             : std_logic;                     -- mm_interconnect_2:Change_Detection_Mem_to_Stream_Translator_master_waitrequest -> Change_Detection_Mem_to_Stream_Translator:master_waitrequest
	signal change_detection_mem_to_stream_translator_master_address                                 : std_logic_vector(1 downto 0);  -- Change_Detection_Mem_to_Stream_Translator:master_address -> mm_interconnect_2:Change_Detection_Mem_to_Stream_Translator_master_address
	signal change_detection_mem_to_stream_translator_master_byteenable                              : std_logic_vector(3 downto 0);  -- Change_Detection_Mem_to_Stream_Translator:master_byteenable -> mm_interconnect_2:Change_Detection_Mem_to_Stream_Translator_master_byteenable
	signal change_detection_mem_to_stream_translator_master_read                                    : std_logic;                     -- Change_Detection_Mem_to_Stream_Translator:master_read -> mm_interconnect_2:Change_Detection_Mem_to_Stream_Translator_master_read
	signal change_detection_mem_to_stream_translator_master_write                                   : std_logic;                     -- Change_Detection_Mem_to_Stream_Translator:master_write -> mm_interconnect_2:Change_Detection_Mem_to_Stream_Translator_master_write
	signal change_detection_mem_to_stream_translator_master_writedata                               : std_logic_vector(31 downto 0); -- Change_Detection_Mem_to_Stream_Translator:master_writedata -> mm_interconnect_2:Change_Detection_Mem_to_Stream_Translator_master_writedata
	signal mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_readdata   : std_logic_vector(31 downto 0); -- Change_Detection_Mem_to_Stream_DMA:slave_readdata -> mm_interconnect_2:Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_readdata
	signal mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_2:Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_address -> Change_Detection_Mem_to_Stream_DMA:slave_address
	signal mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_read       : std_logic;                     -- mm_interconnect_2:Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_read -> Change_Detection_Mem_to_Stream_DMA:slave_read
	signal mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_2:Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_byteenable -> Change_Detection_Mem_to_Stream_DMA:slave_byteenable
	signal mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_write      : std_logic;                     -- mm_interconnect_2:Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_write -> Change_Detection_Mem_to_Stream_DMA:slave_write
	signal mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_2:Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_writedata -> Change_Detection_Mem_to_Stream_DMA:slave_writedata
	signal change_detection_stream_to_mem_translator_master_readdata                                : std_logic_vector(31 downto 0); -- mm_interconnect_3:Change_Detection_Stream_to_Mem_Translator_master_readdata -> Change_Detection_Stream_to_Mem_Translator:master_readdata
	signal change_detection_stream_to_mem_translator_master_waitrequest                             : std_logic;                     -- mm_interconnect_3:Change_Detection_Stream_to_Mem_Translator_master_waitrequest -> Change_Detection_Stream_to_Mem_Translator:master_waitrequest
	signal change_detection_stream_to_mem_translator_master_address                                 : std_logic_vector(1 downto 0);  -- Change_Detection_Stream_to_Mem_Translator:master_address -> mm_interconnect_3:Change_Detection_Stream_to_Mem_Translator_master_address
	signal change_detection_stream_to_mem_translator_master_byteenable                              : std_logic_vector(3 downto 0);  -- Change_Detection_Stream_to_Mem_Translator:master_byteenable -> mm_interconnect_3:Change_Detection_Stream_to_Mem_Translator_master_byteenable
	signal change_detection_stream_to_mem_translator_master_read                                    : std_logic;                     -- Change_Detection_Stream_to_Mem_Translator:master_read -> mm_interconnect_3:Change_Detection_Stream_to_Mem_Translator_master_read
	signal change_detection_stream_to_mem_translator_master_write                                   : std_logic;                     -- Change_Detection_Stream_to_Mem_Translator:master_write -> mm_interconnect_3:Change_Detection_Stream_to_Mem_Translator_master_write
	signal change_detection_stream_to_mem_translator_master_writedata                               : std_logic_vector(31 downto 0); -- Change_Detection_Stream_to_Mem_Translator:master_writedata -> mm_interconnect_3:Change_Detection_Stream_to_Mem_Translator_master_writedata
	signal mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_readdata   : std_logic_vector(31 downto 0); -- Change_Detection_Stream_to_Mem_DMA:slave_readdata -> mm_interconnect_3:Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_readdata
	signal mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_3:Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_address -> Change_Detection_Stream_to_Mem_DMA:slave_address
	signal mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_read       : std_logic;                     -- mm_interconnect_3:Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_read -> Change_Detection_Stream_to_Mem_DMA:slave_read
	signal mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_3:Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_byteenable -> Change_Detection_Stream_to_Mem_DMA:slave_byteenable
	signal mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_write      : std_logic;                     -- mm_interconnect_3:Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_write -> Change_Detection_Stream_to_Mem_DMA:slave_write
	signal mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_3:Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_writedata -> Change_Detection_Stream_to_Mem_DMA:slave_writedata
	signal arm_a9_hps_f2h_irq0_irq                                                                  : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p0
	signal arm_a9_hps_f2h_irq1_irq                                                                  : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	signal rst_controller_reset_out_reset                                                           : std_logic;                     -- rst_controller:reset_out -> [Anomaly_Detection_Module:rst, Change_Detection_Mem_to_Stream_DMA:reset, Change_Detection_Mem_to_Stream_Translator:reset, Change_Detection_Stream_to_Mem_DMA:reset, Change_Detection_Stream_to_Mem_Translator:reset, mm_interconnect_0:Change_Detection_Mem_to_Stream_DMA_reset_reset_bridge_in_reset_reset, mm_interconnect_1:Change_Detection_Mem_to_Stream_Translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:Change_Detection_Mem_to_Stream_Translator_reset_reset_bridge_in_reset_reset, mm_interconnect_3:Change_Detection_Stream_to_Mem_Translator_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal arm_a9_hps_h2f_reset_reset                                                               : std_logic;                     -- ARM_A9_HPS:h2f_rst_n -> arm_a9_hps_h2f_reset_reset:in
	signal system_pll_reset_source_reset                                                            : std_logic;                     -- System_PLL:reset_source_reset -> rst_controller:reset_in1
	signal rst_controller_001_reset_out_reset                                                       : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	signal mm_interconnect_0_sdram_s1_read_ports_inv                                                : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> SDRAM:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> SDRAM:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                                               : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> SDRAM:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                                                 : std_logic;                     -- rst_controller_reset_out_reset:inv -> SDRAM:reset_n
	signal arm_a9_hps_h2f_reset_reset_ports_inv                                                     : std_logic;                     -- arm_a9_hps_h2f_reset_reset:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]

begin

	arm_a9_hps : component dma_platform_ARM_A9_HPS
		generic map (
			F2S_Width => 2,
			S2F_Width => 2
		)
		port map (
			f2h_stm_hwevents         => arm_a9_hps_f2h_stm_hw_events_stm_hwevents, -- f2h_stm_hw_events.stm_hwevents
			mem_a                    => memory_mem_a,                              --            memory.mem_a
			mem_ba                   => memory_mem_ba,                             --                  .mem_ba
			mem_ck                   => memory_mem_ck,                             --                  .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                           --                  .mem_ck_n
			mem_cke                  => memory_mem_cke,                            --                  .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                           --                  .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                          --                  .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                          --                  .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                           --                  .mem_we_n
			mem_reset_n              => memory_mem_reset_n,                        --                  .mem_reset_n
			mem_dq                   => memory_mem_dq,                             --                  .mem_dq
			mem_dqs                  => memory_mem_dqs,                            --                  .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                          --                  .mem_dqs_n
			mem_odt                  => memory_mem_odt,                            --                  .mem_odt
			mem_dm                   => memory_mem_dm,                             --                  .mem_dm
			oct_rzqin                => memory_oct_rzqin,                          --                  .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_io_hps_io_emac1_inst_TX_CLK,           --            hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_io_hps_io_emac1_inst_TXD0,             --                  .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_io_hps_io_emac1_inst_TXD1,             --                  .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_io_hps_io_emac1_inst_TXD2,             --                  .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_io_hps_io_emac1_inst_TXD3,             --                  .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_io_hps_io_emac1_inst_RXD0,             --                  .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_io_hps_io_emac1_inst_MDIO,             --                  .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_io_hps_io_emac1_inst_MDC,              --                  .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_io_hps_io_emac1_inst_RX_CTL,           --                  .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_io_hps_io_emac1_inst_TX_CTL,           --                  .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_io_hps_io_emac1_inst_RX_CLK,           --                  .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_io_hps_io_emac1_inst_RXD1,             --                  .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_io_hps_io_emac1_inst_RXD2,             --                  .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_io_hps_io_emac1_inst_RXD3,             --                  .hps_io_emac1_inst_RXD3
			hps_io_qspi_inst_IO0     => hps_io_hps_io_qspi_inst_IO0,               --                  .hps_io_qspi_inst_IO0
			hps_io_qspi_inst_IO1     => hps_io_hps_io_qspi_inst_IO1,               --                  .hps_io_qspi_inst_IO1
			hps_io_qspi_inst_IO2     => hps_io_hps_io_qspi_inst_IO2,               --                  .hps_io_qspi_inst_IO2
			hps_io_qspi_inst_IO3     => hps_io_hps_io_qspi_inst_IO3,               --                  .hps_io_qspi_inst_IO3
			hps_io_qspi_inst_SS0     => hps_io_hps_io_qspi_inst_SS0,               --                  .hps_io_qspi_inst_SS0
			hps_io_qspi_inst_CLK     => hps_io_hps_io_qspi_inst_CLK,               --                  .hps_io_qspi_inst_CLK
			hps_io_sdio_inst_CMD     => hps_io_hps_io_sdio_inst_CMD,               --                  .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_io_hps_io_sdio_inst_D0,                --                  .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_io_hps_io_sdio_inst_D1,                --                  .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_io_hps_io_sdio_inst_CLK,               --                  .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_io_hps_io_sdio_inst_D2,                --                  .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_io_hps_io_sdio_inst_D3,                --                  .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_io_hps_io_usb1_inst_D0,                --                  .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_io_hps_io_usb1_inst_D1,                --                  .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_io_hps_io_usb1_inst_D2,                --                  .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_io_hps_io_usb1_inst_D3,                --                  .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_io_hps_io_usb1_inst_D4,                --                  .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_io_hps_io_usb1_inst_D5,                --                  .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_io_hps_io_usb1_inst_D6,                --                  .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_io_hps_io_usb1_inst_D7,                --                  .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_io_hps_io_usb1_inst_CLK,               --                  .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_io_hps_io_usb1_inst_STP,               --                  .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_io_hps_io_usb1_inst_DIR,               --                  .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_io_hps_io_usb1_inst_NXT,               --                  .hps_io_usb1_inst_NXT
			hps_io_spim0_inst_CLK    => hps_io_hps_io_spim0_inst_CLK,              --                  .hps_io_spim0_inst_CLK
			hps_io_spim0_inst_MOSI   => hps_io_hps_io_spim0_inst_MOSI,             --                  .hps_io_spim0_inst_MOSI
			hps_io_spim0_inst_MISO   => hps_io_hps_io_spim0_inst_MISO,             --                  .hps_io_spim0_inst_MISO
			hps_io_spim0_inst_SS0    => hps_io_hps_io_spim0_inst_SS0,              --                  .hps_io_spim0_inst_SS0
			hps_io_spim1_inst_CLK    => hps_io_hps_io_spim1_inst_CLK,              --                  .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   => hps_io_hps_io_spim1_inst_MOSI,             --                  .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   => hps_io_hps_io_spim1_inst_MISO,             --                  .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    => hps_io_hps_io_spim1_inst_SS0,              --                  .hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     => hps_io_hps_io_uart0_inst_RX,               --                  .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_io_hps_io_uart0_inst_TX,               --                  .hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     => hps_io_hps_io_i2c0_inst_SDA,               --                  .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     => hps_io_hps_io_i2c0_inst_SCL,               --                  .hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     => hps_io_hps_io_i2c1_inst_SDA,               --                  .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_io_hps_io_i2c1_inst_SCL,               --                  .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  => hps_io_hps_io_gpio_inst_GPIO09,            --                  .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  => hps_io_hps_io_gpio_inst_GPIO35,            --                  .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO37  => hps_io_hps_io_gpio_inst_GPIO37,            --                  .hps_io_gpio_inst_GPIO37
			hps_io_gpio_inst_GPIO40  => hps_io_hps_io_gpio_inst_GPIO40,            --                  .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO41  => hps_io_hps_io_gpio_inst_GPIO41,            --                  .hps_io_gpio_inst_GPIO41
			hps_io_gpio_inst_GPIO44  => hps_io_hps_io_gpio_inst_GPIO44,            --                  .hps_io_gpio_inst_GPIO44
			hps_io_gpio_inst_GPIO48  => hps_io_hps_io_gpio_inst_GPIO48,            --                  .hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  => hps_io_hps_io_gpio_inst_GPIO53,            --                  .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_io_hps_io_gpio_inst_GPIO54,            --                  .hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  => hps_io_hps_io_gpio_inst_GPIO61,            --                  .hps_io_gpio_inst_GPIO61
			h2f_rst_n                => arm_a9_hps_h2f_reset_reset,                --         h2f_reset.reset_n
			h2f_axi_clk              => system_pll_sys_clk_clk,                    --     h2f_axi_clock.clk
			h2f_AWID                 => arm_a9_hps_h2f_axi_master_awid,            --    h2f_axi_master.awid
			h2f_AWADDR               => arm_a9_hps_h2f_axi_master_awaddr,          --                  .awaddr
			h2f_AWLEN                => arm_a9_hps_h2f_axi_master_awlen,           --                  .awlen
			h2f_AWSIZE               => arm_a9_hps_h2f_axi_master_awsize,          --                  .awsize
			h2f_AWBURST              => arm_a9_hps_h2f_axi_master_awburst,         --                  .awburst
			h2f_AWLOCK               => arm_a9_hps_h2f_axi_master_awlock,          --                  .awlock
			h2f_AWCACHE              => arm_a9_hps_h2f_axi_master_awcache,         --                  .awcache
			h2f_AWPROT               => arm_a9_hps_h2f_axi_master_awprot,          --                  .awprot
			h2f_AWVALID              => arm_a9_hps_h2f_axi_master_awvalid,         --                  .awvalid
			h2f_AWREADY              => arm_a9_hps_h2f_axi_master_awready,         --                  .awready
			h2f_WID                  => arm_a9_hps_h2f_axi_master_wid,             --                  .wid
			h2f_WDATA                => arm_a9_hps_h2f_axi_master_wdata,           --                  .wdata
			h2f_WSTRB                => arm_a9_hps_h2f_axi_master_wstrb,           --                  .wstrb
			h2f_WLAST                => arm_a9_hps_h2f_axi_master_wlast,           --                  .wlast
			h2f_WVALID               => arm_a9_hps_h2f_axi_master_wvalid,          --                  .wvalid
			h2f_WREADY               => arm_a9_hps_h2f_axi_master_wready,          --                  .wready
			h2f_BID                  => arm_a9_hps_h2f_axi_master_bid,             --                  .bid
			h2f_BRESP                => arm_a9_hps_h2f_axi_master_bresp,           --                  .bresp
			h2f_BVALID               => arm_a9_hps_h2f_axi_master_bvalid,          --                  .bvalid
			h2f_BREADY               => arm_a9_hps_h2f_axi_master_bready,          --                  .bready
			h2f_ARID                 => arm_a9_hps_h2f_axi_master_arid,            --                  .arid
			h2f_ARADDR               => arm_a9_hps_h2f_axi_master_araddr,          --                  .araddr
			h2f_ARLEN                => arm_a9_hps_h2f_axi_master_arlen,           --                  .arlen
			h2f_ARSIZE               => arm_a9_hps_h2f_axi_master_arsize,          --                  .arsize
			h2f_ARBURST              => arm_a9_hps_h2f_axi_master_arburst,         --                  .arburst
			h2f_ARLOCK               => arm_a9_hps_h2f_axi_master_arlock,          --                  .arlock
			h2f_ARCACHE              => arm_a9_hps_h2f_axi_master_arcache,         --                  .arcache
			h2f_ARPROT               => arm_a9_hps_h2f_axi_master_arprot,          --                  .arprot
			h2f_ARVALID              => arm_a9_hps_h2f_axi_master_arvalid,         --                  .arvalid
			h2f_ARREADY              => arm_a9_hps_h2f_axi_master_arready,         --                  .arready
			h2f_RID                  => arm_a9_hps_h2f_axi_master_rid,             --                  .rid
			h2f_RDATA                => arm_a9_hps_h2f_axi_master_rdata,           --                  .rdata
			h2f_RRESP                => arm_a9_hps_h2f_axi_master_rresp,           --                  .rresp
			h2f_RLAST                => arm_a9_hps_h2f_axi_master_rlast,           --                  .rlast
			h2f_RVALID               => arm_a9_hps_h2f_axi_master_rvalid,          --                  .rvalid
			h2f_RREADY               => arm_a9_hps_h2f_axi_master_rready,          --                  .rready
			f2h_axi_clk              => system_pll_sys_clk_clk,                    --     f2h_axi_clock.clk
			f2h_AWID                 => open,                                      --     f2h_axi_slave.awid
			f2h_AWADDR               => open,                                      --                  .awaddr
			f2h_AWLEN                => open,                                      --                  .awlen
			f2h_AWSIZE               => open,                                      --                  .awsize
			f2h_AWBURST              => open,                                      --                  .awburst
			f2h_AWLOCK               => open,                                      --                  .awlock
			f2h_AWCACHE              => open,                                      --                  .awcache
			f2h_AWPROT               => open,                                      --                  .awprot
			f2h_AWVALID              => open,                                      --                  .awvalid
			f2h_AWREADY              => open,                                      --                  .awready
			f2h_AWUSER               => open,                                      --                  .awuser
			f2h_WID                  => open,                                      --                  .wid
			f2h_WDATA                => open,                                      --                  .wdata
			f2h_WSTRB                => open,                                      --                  .wstrb
			f2h_WLAST                => open,                                      --                  .wlast
			f2h_WVALID               => open,                                      --                  .wvalid
			f2h_WREADY               => open,                                      --                  .wready
			f2h_BID                  => open,                                      --                  .bid
			f2h_BRESP                => open,                                      --                  .bresp
			f2h_BVALID               => open,                                      --                  .bvalid
			f2h_BREADY               => open,                                      --                  .bready
			f2h_ARID                 => open,                                      --                  .arid
			f2h_ARADDR               => open,                                      --                  .araddr
			f2h_ARLEN                => open,                                      --                  .arlen
			f2h_ARSIZE               => open,                                      --                  .arsize
			f2h_ARBURST              => open,                                      --                  .arburst
			f2h_ARLOCK               => open,                                      --                  .arlock
			f2h_ARCACHE              => open,                                      --                  .arcache
			f2h_ARPROT               => open,                                      --                  .arprot
			f2h_ARVALID              => open,                                      --                  .arvalid
			f2h_ARREADY              => open,                                      --                  .arready
			f2h_ARUSER               => open,                                      --                  .aruser
			f2h_RID                  => open,                                      --                  .rid
			f2h_RDATA                => open,                                      --                  .rdata
			f2h_RRESP                => open,                                      --                  .rresp
			f2h_RLAST                => open,                                      --                  .rlast
			f2h_RVALID               => open,                                      --                  .rvalid
			f2h_RREADY               => open,                                      --                  .rready
			h2f_lw_axi_clk           => system_pll_sys_clk_clk,                    --  h2f_lw_axi_clock.clk
			h2f_lw_AWID              => arm_a9_hps_h2f_lw_axi_master_awid,         -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => arm_a9_hps_h2f_lw_axi_master_awaddr,       --                  .awaddr
			h2f_lw_AWLEN             => arm_a9_hps_h2f_lw_axi_master_awlen,        --                  .awlen
			h2f_lw_AWSIZE            => arm_a9_hps_h2f_lw_axi_master_awsize,       --                  .awsize
			h2f_lw_AWBURST           => arm_a9_hps_h2f_lw_axi_master_awburst,      --                  .awburst
			h2f_lw_AWLOCK            => arm_a9_hps_h2f_lw_axi_master_awlock,       --                  .awlock
			h2f_lw_AWCACHE           => arm_a9_hps_h2f_lw_axi_master_awcache,      --                  .awcache
			h2f_lw_AWPROT            => arm_a9_hps_h2f_lw_axi_master_awprot,       --                  .awprot
			h2f_lw_AWVALID           => arm_a9_hps_h2f_lw_axi_master_awvalid,      --                  .awvalid
			h2f_lw_AWREADY           => arm_a9_hps_h2f_lw_axi_master_awready,      --                  .awready
			h2f_lw_WID               => arm_a9_hps_h2f_lw_axi_master_wid,          --                  .wid
			h2f_lw_WDATA             => arm_a9_hps_h2f_lw_axi_master_wdata,        --                  .wdata
			h2f_lw_WSTRB             => arm_a9_hps_h2f_lw_axi_master_wstrb,        --                  .wstrb
			h2f_lw_WLAST             => arm_a9_hps_h2f_lw_axi_master_wlast,        --                  .wlast
			h2f_lw_WVALID            => arm_a9_hps_h2f_lw_axi_master_wvalid,       --                  .wvalid
			h2f_lw_WREADY            => arm_a9_hps_h2f_lw_axi_master_wready,       --                  .wready
			h2f_lw_BID               => arm_a9_hps_h2f_lw_axi_master_bid,          --                  .bid
			h2f_lw_BRESP             => arm_a9_hps_h2f_lw_axi_master_bresp,        --                  .bresp
			h2f_lw_BVALID            => arm_a9_hps_h2f_lw_axi_master_bvalid,       --                  .bvalid
			h2f_lw_BREADY            => arm_a9_hps_h2f_lw_axi_master_bready,       --                  .bready
			h2f_lw_ARID              => arm_a9_hps_h2f_lw_axi_master_arid,         --                  .arid
			h2f_lw_ARADDR            => arm_a9_hps_h2f_lw_axi_master_araddr,       --                  .araddr
			h2f_lw_ARLEN             => arm_a9_hps_h2f_lw_axi_master_arlen,        --                  .arlen
			h2f_lw_ARSIZE            => arm_a9_hps_h2f_lw_axi_master_arsize,       --                  .arsize
			h2f_lw_ARBURST           => arm_a9_hps_h2f_lw_axi_master_arburst,      --                  .arburst
			h2f_lw_ARLOCK            => arm_a9_hps_h2f_lw_axi_master_arlock,       --                  .arlock
			h2f_lw_ARCACHE           => arm_a9_hps_h2f_lw_axi_master_arcache,      --                  .arcache
			h2f_lw_ARPROT            => arm_a9_hps_h2f_lw_axi_master_arprot,       --                  .arprot
			h2f_lw_ARVALID           => arm_a9_hps_h2f_lw_axi_master_arvalid,      --                  .arvalid
			h2f_lw_ARREADY           => arm_a9_hps_h2f_lw_axi_master_arready,      --                  .arready
			h2f_lw_RID               => arm_a9_hps_h2f_lw_axi_master_rid,          --                  .rid
			h2f_lw_RDATA             => arm_a9_hps_h2f_lw_axi_master_rdata,        --                  .rdata
			h2f_lw_RRESP             => arm_a9_hps_h2f_lw_axi_master_rresp,        --                  .rresp
			h2f_lw_RLAST             => arm_a9_hps_h2f_lw_axi_master_rlast,        --                  .rlast
			h2f_lw_RVALID            => arm_a9_hps_h2f_lw_axi_master_rvalid,       --                  .rvalid
			h2f_lw_RREADY            => arm_a9_hps_h2f_lw_axi_master_rready,       --                  .rready
			f2h_irq_p0               => arm_a9_hps_f2h_irq0_irq,                   --          f2h_irq0.irq
			f2h_irq_p1               => arm_a9_hps_f2h_irq1_irq                    --          f2h_irq1.irq
		);

	anomaly_detection_module : component anomaly_detection
		generic map (
			IM_SIZE     => 500,
			ADDR_SIZE   => 16,
			WORD_SIZE   => 16,
			COUNT_WIDTH => 9
		)
		port map (
			clk             => system_pll_sys_clk_clk,                                               --              clock_sink.clk
			rst             => rst_controller_reset_out_reset,                                       --             clock_reset.reset
			data_out        => anomaly_detection_module_avalon_streaming_source_data,                -- avalon_streaming_source.data
			endpacket_out   => anomaly_detection_module_avalon_streaming_source_endofpacket,         --                        .endofpacket
			ready_in        => anomaly_detection_module_avalon_streaming_source_ready,               --                        .ready
			startpacket_out => anomaly_detection_module_avalon_streaming_source_startofpacket,       --                        .startofpacket
			valid_out       => anomaly_detection_module_avalon_streaming_source_valid,               --                        .valid
			data_in         => change_detection_mem_to_stream_dma_avalon_pixel_source_data,          --   avalon_streaming_sink.data
			endpacket_in    => change_detection_mem_to_stream_dma_avalon_pixel_source_endofpacket,   --                        .endofpacket
			ready_out       => change_detection_mem_to_stream_dma_avalon_pixel_source_ready,         --                        .ready
			startpacket_in  => change_detection_mem_to_stream_dma_avalon_pixel_source_startofpacket, --                        .startofpacket
			valid_in        => change_detection_mem_to_stream_dma_avalon_pixel_source_valid          --                        .valid
		);

	change_detection_mem_to_stream_dma : component dma_platform_Change_Detection_Mem_to_Stream_DMA
		port map (
			clk                  => system_pll_sys_clk_clk,                                                                   --                      clk.clk
			reset                => rst_controller_reset_out_reset,                                                           --                    reset.reset
			master_address       => change_detection_mem_to_stream_dma_avalon_dma_master_address,                             --        avalon_dma_master.address
			master_waitrequest   => change_detection_mem_to_stream_dma_avalon_dma_master_waitrequest,                         --                         .waitrequest
			master_arbiterlock   => change_detection_mem_to_stream_dma_avalon_dma_master_lock,                                --                         .lock
			master_read          => change_detection_mem_to_stream_dma_avalon_dma_master_read,                                --                         .read
			master_readdata      => change_detection_mem_to_stream_dma_avalon_dma_master_readdata,                            --                         .readdata
			master_readdatavalid => change_detection_mem_to_stream_dma_avalon_dma_master_readdatavalid,                       --                         .readdatavalid
			slave_address        => mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_address,    -- avalon_dma_control_slave.address
			slave_byteenable     => mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_byteenable, --                         .byteenable
			slave_read           => mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_read,       --                         .read
			slave_write          => mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_write,      --                         .write
			slave_writedata      => mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_writedata,  --                         .writedata
			slave_readdata       => mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_readdata,   --                         .readdata
			stream_ready         => change_detection_mem_to_stream_dma_avalon_pixel_source_ready,                             --      avalon_pixel_source.ready
			stream_data          => change_detection_mem_to_stream_dma_avalon_pixel_source_data,                              --                         .data
			stream_startofpacket => change_detection_mem_to_stream_dma_avalon_pixel_source_startofpacket,                     --                         .startofpacket
			stream_endofpacket   => change_detection_mem_to_stream_dma_avalon_pixel_source_endofpacket,                       --                         .endofpacket
			stream_valid         => change_detection_mem_to_stream_dma_avalon_pixel_source_valid                              --                         .valid
		);

	change_detection_mem_to_stream_translator : component altera_up_avalon_video_dma_ctrl_addr_trans
		generic map (
			ADDRESS_TRANSLATION_MASK => "11000000000000000000000000000000"
		)
		port map (
			clk                => system_pll_sys_clk_clk,                                                        --  clock.clk
			reset              => rst_controller_reset_out_reset,                                                --  reset.reset
			slave_address      => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_address,     --  slave.address
			slave_byteenable   => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_byteenable,  --       .byteenable
			slave_read         => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_read,        --       .read
			slave_write        => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_write,       --       .write
			slave_writedata    => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_writedata,   --       .writedata
			slave_readdata     => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_readdata,    --       .readdata
			slave_waitrequest  => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_waitrequest, --       .waitrequest
			master_readdata    => change_detection_mem_to_stream_translator_master_readdata,                     -- master.readdata
			master_waitrequest => change_detection_mem_to_stream_translator_master_waitrequest,                  --       .waitrequest
			master_address     => change_detection_mem_to_stream_translator_master_address,                      --       .address
			master_byteenable  => change_detection_mem_to_stream_translator_master_byteenable,                   --       .byteenable
			master_read        => change_detection_mem_to_stream_translator_master_read,                         --       .read
			master_write       => change_detection_mem_to_stream_translator_master_write,                        --       .write
			master_writedata   => change_detection_mem_to_stream_translator_master_writedata                     --       .writedata
		);

	change_detection_stream_to_mem_dma : component dma_platform_Change_Detection_Stream_to_Mem_DMA
		port map (
			clk                  => system_pll_sys_clk_clk,                                                                   --                      clk.clk
			reset                => rst_controller_reset_out_reset,                                                           --                    reset.reset
			stream_data          => anomaly_detection_module_avalon_streaming_source_data,                                    --          avalon_dma_sink.data
			stream_startofpacket => anomaly_detection_module_avalon_streaming_source_startofpacket,                           --                         .startofpacket
			stream_endofpacket   => anomaly_detection_module_avalon_streaming_source_endofpacket,                             --                         .endofpacket
			stream_valid         => anomaly_detection_module_avalon_streaming_source_valid,                                   --                         .valid
			stream_ready         => anomaly_detection_module_avalon_streaming_source_ready,                                   --                         .ready
			slave_address        => mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_address,    -- avalon_dma_control_slave.address
			slave_byteenable     => mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_byteenable, --                         .byteenable
			slave_read           => mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_read,       --                         .read
			slave_write          => mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_write,      --                         .write
			slave_writedata      => mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_writedata,  --                         .writedata
			slave_readdata       => mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_readdata,   --                         .readdata
			master_address       => change_detection_stream_to_mem_dma_avalon_dma_master_address,                             --        avalon_dma_master.address
			master_waitrequest   => change_detection_stream_to_mem_dma_avalon_dma_master_waitrequest,                         --                         .waitrequest
			master_write         => change_detection_stream_to_mem_dma_avalon_dma_master_write,                               --                         .write
			master_writedata     => change_detection_stream_to_mem_dma_avalon_dma_master_writedata                            --                         .writedata
		);

	change_detection_stream_to_mem_translator : component altera_up_avalon_video_dma_ctrl_addr_trans
		generic map (
			ADDRESS_TRANSLATION_MASK => "11000000000000000000000000000000"
		)
		port map (
			clk                => system_pll_sys_clk_clk,                                                        --  clock.clk
			reset              => rst_controller_reset_out_reset,                                                --  reset.reset
			slave_address      => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_address,     --  slave.address
			slave_byteenable   => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_byteenable,  --       .byteenable
			slave_read         => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_read,        --       .read
			slave_write        => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_write,       --       .write
			slave_writedata    => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_writedata,   --       .writedata
			slave_readdata     => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_readdata,    --       .readdata
			slave_waitrequest  => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_waitrequest, --       .waitrequest
			master_readdata    => change_detection_stream_to_mem_translator_master_readdata,                     -- master.readdata
			master_waitrequest => change_detection_stream_to_mem_translator_master_waitrequest,                  --       .waitrequest
			master_address     => change_detection_stream_to_mem_translator_master_address,                      --       .address
			master_byteenable  => change_detection_stream_to_mem_translator_master_byteenable,                   --       .byteenable
			master_read        => change_detection_stream_to_mem_translator_master_read,                         --       .read
			master_write       => change_detection_stream_to_mem_translator_master_write,                        --       .write
			master_writedata   => change_detection_stream_to_mem_translator_master_writedata                     --       .writedata
		);

	sdram : component dma_platform_SDRAM
		port map (
			clk            => system_pll_sys_clk_clk,                          --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	system_pll : component dma_platform_System_PLL
		port map (
			ref_clk_clk        => system_pll_ref_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => system_pll_ref_reset_reset,    --    ref_reset.reset
			sys_clk_clk        => system_pll_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => open,                          --    sdram_clk.clk
			reset_source_reset => system_pll_reset_source_reset  -- reset_source.reset
		);

	mm_interconnect_0 : component dma_platform_mm_interconnect_0
		port map (
			ARM_A9_HPS_h2f_axi_master_awid                                        => arm_a9_hps_h2f_axi_master_awid,                                     --                                       ARM_A9_HPS_h2f_axi_master.awid
			ARM_A9_HPS_h2f_axi_master_awaddr                                      => arm_a9_hps_h2f_axi_master_awaddr,                                   --                                                                .awaddr
			ARM_A9_HPS_h2f_axi_master_awlen                                       => arm_a9_hps_h2f_axi_master_awlen,                                    --                                                                .awlen
			ARM_A9_HPS_h2f_axi_master_awsize                                      => arm_a9_hps_h2f_axi_master_awsize,                                   --                                                                .awsize
			ARM_A9_HPS_h2f_axi_master_awburst                                     => arm_a9_hps_h2f_axi_master_awburst,                                  --                                                                .awburst
			ARM_A9_HPS_h2f_axi_master_awlock                                      => arm_a9_hps_h2f_axi_master_awlock,                                   --                                                                .awlock
			ARM_A9_HPS_h2f_axi_master_awcache                                     => arm_a9_hps_h2f_axi_master_awcache,                                  --                                                                .awcache
			ARM_A9_HPS_h2f_axi_master_awprot                                      => arm_a9_hps_h2f_axi_master_awprot,                                   --                                                                .awprot
			ARM_A9_HPS_h2f_axi_master_awvalid                                     => arm_a9_hps_h2f_axi_master_awvalid,                                  --                                                                .awvalid
			ARM_A9_HPS_h2f_axi_master_awready                                     => arm_a9_hps_h2f_axi_master_awready,                                  --                                                                .awready
			ARM_A9_HPS_h2f_axi_master_wid                                         => arm_a9_hps_h2f_axi_master_wid,                                      --                                                                .wid
			ARM_A9_HPS_h2f_axi_master_wdata                                       => arm_a9_hps_h2f_axi_master_wdata,                                    --                                                                .wdata
			ARM_A9_HPS_h2f_axi_master_wstrb                                       => arm_a9_hps_h2f_axi_master_wstrb,                                    --                                                                .wstrb
			ARM_A9_HPS_h2f_axi_master_wlast                                       => arm_a9_hps_h2f_axi_master_wlast,                                    --                                                                .wlast
			ARM_A9_HPS_h2f_axi_master_wvalid                                      => arm_a9_hps_h2f_axi_master_wvalid,                                   --                                                                .wvalid
			ARM_A9_HPS_h2f_axi_master_wready                                      => arm_a9_hps_h2f_axi_master_wready,                                   --                                                                .wready
			ARM_A9_HPS_h2f_axi_master_bid                                         => arm_a9_hps_h2f_axi_master_bid,                                      --                                                                .bid
			ARM_A9_HPS_h2f_axi_master_bresp                                       => arm_a9_hps_h2f_axi_master_bresp,                                    --                                                                .bresp
			ARM_A9_HPS_h2f_axi_master_bvalid                                      => arm_a9_hps_h2f_axi_master_bvalid,                                   --                                                                .bvalid
			ARM_A9_HPS_h2f_axi_master_bready                                      => arm_a9_hps_h2f_axi_master_bready,                                   --                                                                .bready
			ARM_A9_HPS_h2f_axi_master_arid                                        => arm_a9_hps_h2f_axi_master_arid,                                     --                                                                .arid
			ARM_A9_HPS_h2f_axi_master_araddr                                      => arm_a9_hps_h2f_axi_master_araddr,                                   --                                                                .araddr
			ARM_A9_HPS_h2f_axi_master_arlen                                       => arm_a9_hps_h2f_axi_master_arlen,                                    --                                                                .arlen
			ARM_A9_HPS_h2f_axi_master_arsize                                      => arm_a9_hps_h2f_axi_master_arsize,                                   --                                                                .arsize
			ARM_A9_HPS_h2f_axi_master_arburst                                     => arm_a9_hps_h2f_axi_master_arburst,                                  --                                                                .arburst
			ARM_A9_HPS_h2f_axi_master_arlock                                      => arm_a9_hps_h2f_axi_master_arlock,                                   --                                                                .arlock
			ARM_A9_HPS_h2f_axi_master_arcache                                     => arm_a9_hps_h2f_axi_master_arcache,                                  --                                                                .arcache
			ARM_A9_HPS_h2f_axi_master_arprot                                      => arm_a9_hps_h2f_axi_master_arprot,                                   --                                                                .arprot
			ARM_A9_HPS_h2f_axi_master_arvalid                                     => arm_a9_hps_h2f_axi_master_arvalid,                                  --                                                                .arvalid
			ARM_A9_HPS_h2f_axi_master_arready                                     => arm_a9_hps_h2f_axi_master_arready,                                  --                                                                .arready
			ARM_A9_HPS_h2f_axi_master_rid                                         => arm_a9_hps_h2f_axi_master_rid,                                      --                                                                .rid
			ARM_A9_HPS_h2f_axi_master_rdata                                       => arm_a9_hps_h2f_axi_master_rdata,                                    --                                                                .rdata
			ARM_A9_HPS_h2f_axi_master_rresp                                       => arm_a9_hps_h2f_axi_master_rresp,                                    --                                                                .rresp
			ARM_A9_HPS_h2f_axi_master_rlast                                       => arm_a9_hps_h2f_axi_master_rlast,                                    --                                                                .rlast
			ARM_A9_HPS_h2f_axi_master_rvalid                                      => arm_a9_hps_h2f_axi_master_rvalid,                                   --                                                                .rvalid
			ARM_A9_HPS_h2f_axi_master_rready                                      => arm_a9_hps_h2f_axi_master_rready,                                   --                                                                .rready
			System_PLL_sys_clk_clk                                                => system_pll_sys_clk_clk,                                             --                                              System_PLL_sys_clk.clk
			ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                                 -- ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			Change_Detection_Mem_to_Stream_DMA_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                                     --  Change_Detection_Mem_to_Stream_DMA_reset_reset_bridge_in_reset.reset
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_address          => change_detection_mem_to_stream_dma_avalon_dma_master_address,       --            Change_Detection_Mem_to_Stream_DMA_avalon_dma_master.address
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_waitrequest      => change_detection_mem_to_stream_dma_avalon_dma_master_waitrequest,   --                                                                .waitrequest
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_read             => change_detection_mem_to_stream_dma_avalon_dma_master_read,          --                                                                .read
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_readdata         => change_detection_mem_to_stream_dma_avalon_dma_master_readdata,      --                                                                .readdata
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_readdatavalid    => change_detection_mem_to_stream_dma_avalon_dma_master_readdatavalid, --                                                                .readdatavalid
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_master_lock             => change_detection_mem_to_stream_dma_avalon_dma_master_lock,          --                                                                .lock
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_master_address          => change_detection_stream_to_mem_dma_avalon_dma_master_address,       --            Change_Detection_Stream_to_Mem_DMA_avalon_dma_master.address
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_master_waitrequest      => change_detection_stream_to_mem_dma_avalon_dma_master_waitrequest,   --                                                                .waitrequest
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_master_write            => change_detection_stream_to_mem_dma_avalon_dma_master_write,         --                                                                .write
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_master_writedata        => change_detection_stream_to_mem_dma_avalon_dma_master_writedata,     --                                                                .writedata
			SDRAM_s1_address                                                      => mm_interconnect_0_sdram_s1_address,                                 --                                                        SDRAM_s1.address
			SDRAM_s1_write                                                        => mm_interconnect_0_sdram_s1_write,                                   --                                                                .write
			SDRAM_s1_read                                                         => mm_interconnect_0_sdram_s1_read,                                    --                                                                .read
			SDRAM_s1_readdata                                                     => mm_interconnect_0_sdram_s1_readdata,                                --                                                                .readdata
			SDRAM_s1_writedata                                                    => mm_interconnect_0_sdram_s1_writedata,                               --                                                                .writedata
			SDRAM_s1_byteenable                                                   => mm_interconnect_0_sdram_s1_byteenable,                              --                                                                .byteenable
			SDRAM_s1_readdatavalid                                                => mm_interconnect_0_sdram_s1_readdatavalid,                           --                                                                .readdatavalid
			SDRAM_s1_waitrequest                                                  => mm_interconnect_0_sdram_s1_waitrequest,                             --                                                                .waitrequest
			SDRAM_s1_chipselect                                                   => mm_interconnect_0_sdram_s1_chipselect                               --                                                                .chipselect
		);

	mm_interconnect_1 : component dma_platform_mm_interconnect_1
		port map (
			ARM_A9_HPS_h2f_lw_axi_master_awid                                           => arm_a9_hps_h2f_lw_axi_master_awid,                                             --                                          ARM_A9_HPS_h2f_lw_axi_master.awid
			ARM_A9_HPS_h2f_lw_axi_master_awaddr                                         => arm_a9_hps_h2f_lw_axi_master_awaddr,                                           --                                                                      .awaddr
			ARM_A9_HPS_h2f_lw_axi_master_awlen                                          => arm_a9_hps_h2f_lw_axi_master_awlen,                                            --                                                                      .awlen
			ARM_A9_HPS_h2f_lw_axi_master_awsize                                         => arm_a9_hps_h2f_lw_axi_master_awsize,                                           --                                                                      .awsize
			ARM_A9_HPS_h2f_lw_axi_master_awburst                                        => arm_a9_hps_h2f_lw_axi_master_awburst,                                          --                                                                      .awburst
			ARM_A9_HPS_h2f_lw_axi_master_awlock                                         => arm_a9_hps_h2f_lw_axi_master_awlock,                                           --                                                                      .awlock
			ARM_A9_HPS_h2f_lw_axi_master_awcache                                        => arm_a9_hps_h2f_lw_axi_master_awcache,                                          --                                                                      .awcache
			ARM_A9_HPS_h2f_lw_axi_master_awprot                                         => arm_a9_hps_h2f_lw_axi_master_awprot,                                           --                                                                      .awprot
			ARM_A9_HPS_h2f_lw_axi_master_awvalid                                        => arm_a9_hps_h2f_lw_axi_master_awvalid,                                          --                                                                      .awvalid
			ARM_A9_HPS_h2f_lw_axi_master_awready                                        => arm_a9_hps_h2f_lw_axi_master_awready,                                          --                                                                      .awready
			ARM_A9_HPS_h2f_lw_axi_master_wid                                            => arm_a9_hps_h2f_lw_axi_master_wid,                                              --                                                                      .wid
			ARM_A9_HPS_h2f_lw_axi_master_wdata                                          => arm_a9_hps_h2f_lw_axi_master_wdata,                                            --                                                                      .wdata
			ARM_A9_HPS_h2f_lw_axi_master_wstrb                                          => arm_a9_hps_h2f_lw_axi_master_wstrb,                                            --                                                                      .wstrb
			ARM_A9_HPS_h2f_lw_axi_master_wlast                                          => arm_a9_hps_h2f_lw_axi_master_wlast,                                            --                                                                      .wlast
			ARM_A9_HPS_h2f_lw_axi_master_wvalid                                         => arm_a9_hps_h2f_lw_axi_master_wvalid,                                           --                                                                      .wvalid
			ARM_A9_HPS_h2f_lw_axi_master_wready                                         => arm_a9_hps_h2f_lw_axi_master_wready,                                           --                                                                      .wready
			ARM_A9_HPS_h2f_lw_axi_master_bid                                            => arm_a9_hps_h2f_lw_axi_master_bid,                                              --                                                                      .bid
			ARM_A9_HPS_h2f_lw_axi_master_bresp                                          => arm_a9_hps_h2f_lw_axi_master_bresp,                                            --                                                                      .bresp
			ARM_A9_HPS_h2f_lw_axi_master_bvalid                                         => arm_a9_hps_h2f_lw_axi_master_bvalid,                                           --                                                                      .bvalid
			ARM_A9_HPS_h2f_lw_axi_master_bready                                         => arm_a9_hps_h2f_lw_axi_master_bready,                                           --                                                                      .bready
			ARM_A9_HPS_h2f_lw_axi_master_arid                                           => arm_a9_hps_h2f_lw_axi_master_arid,                                             --                                                                      .arid
			ARM_A9_HPS_h2f_lw_axi_master_araddr                                         => arm_a9_hps_h2f_lw_axi_master_araddr,                                           --                                                                      .araddr
			ARM_A9_HPS_h2f_lw_axi_master_arlen                                          => arm_a9_hps_h2f_lw_axi_master_arlen,                                            --                                                                      .arlen
			ARM_A9_HPS_h2f_lw_axi_master_arsize                                         => arm_a9_hps_h2f_lw_axi_master_arsize,                                           --                                                                      .arsize
			ARM_A9_HPS_h2f_lw_axi_master_arburst                                        => arm_a9_hps_h2f_lw_axi_master_arburst,                                          --                                                                      .arburst
			ARM_A9_HPS_h2f_lw_axi_master_arlock                                         => arm_a9_hps_h2f_lw_axi_master_arlock,                                           --                                                                      .arlock
			ARM_A9_HPS_h2f_lw_axi_master_arcache                                        => arm_a9_hps_h2f_lw_axi_master_arcache,                                          --                                                                      .arcache
			ARM_A9_HPS_h2f_lw_axi_master_arprot                                         => arm_a9_hps_h2f_lw_axi_master_arprot,                                           --                                                                      .arprot
			ARM_A9_HPS_h2f_lw_axi_master_arvalid                                        => arm_a9_hps_h2f_lw_axi_master_arvalid,                                          --                                                                      .arvalid
			ARM_A9_HPS_h2f_lw_axi_master_arready                                        => arm_a9_hps_h2f_lw_axi_master_arready,                                          --                                                                      .arready
			ARM_A9_HPS_h2f_lw_axi_master_rid                                            => arm_a9_hps_h2f_lw_axi_master_rid,                                              --                                                                      .rid
			ARM_A9_HPS_h2f_lw_axi_master_rdata                                          => arm_a9_hps_h2f_lw_axi_master_rdata,                                            --                                                                      .rdata
			ARM_A9_HPS_h2f_lw_axi_master_rresp                                          => arm_a9_hps_h2f_lw_axi_master_rresp,                                            --                                                                      .rresp
			ARM_A9_HPS_h2f_lw_axi_master_rlast                                          => arm_a9_hps_h2f_lw_axi_master_rlast,                                            --                                                                      .rlast
			ARM_A9_HPS_h2f_lw_axi_master_rvalid                                         => arm_a9_hps_h2f_lw_axi_master_rvalid,                                           --                                                                      .rvalid
			ARM_A9_HPS_h2f_lw_axi_master_rready                                         => arm_a9_hps_h2f_lw_axi_master_rready,                                           --                                                                      .rready
			System_PLL_sys_clk_clk                                                      => system_pll_sys_clk_clk,                                                        --                                                    System_PLL_sys_clk.clk
			ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset    => rst_controller_001_reset_out_reset,                                            --    ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			Change_Detection_Mem_to_Stream_Translator_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                                -- Change_Detection_Mem_to_Stream_Translator_reset_reset_bridge_in_reset.reset
			Change_Detection_Mem_to_Stream_Translator_slave_address                     => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_address,     --                       Change_Detection_Mem_to_Stream_Translator_slave.address
			Change_Detection_Mem_to_Stream_Translator_slave_write                       => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_write,       --                                                                      .write
			Change_Detection_Mem_to_Stream_Translator_slave_read                        => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_read,        --                                                                      .read
			Change_Detection_Mem_to_Stream_Translator_slave_readdata                    => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_readdata,    --                                                                      .readdata
			Change_Detection_Mem_to_Stream_Translator_slave_writedata                   => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_writedata,   --                                                                      .writedata
			Change_Detection_Mem_to_Stream_Translator_slave_byteenable                  => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_byteenable,  --                                                                      .byteenable
			Change_Detection_Mem_to_Stream_Translator_slave_waitrequest                 => mm_interconnect_1_change_detection_mem_to_stream_translator_slave_waitrequest, --                                                                      .waitrequest
			Change_Detection_Stream_to_Mem_Translator_slave_address                     => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_address,     --                       Change_Detection_Stream_to_Mem_Translator_slave.address
			Change_Detection_Stream_to_Mem_Translator_slave_write                       => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_write,       --                                                                      .write
			Change_Detection_Stream_to_Mem_Translator_slave_read                        => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_read,        --                                                                      .read
			Change_Detection_Stream_to_Mem_Translator_slave_readdata                    => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_readdata,    --                                                                      .readdata
			Change_Detection_Stream_to_Mem_Translator_slave_writedata                   => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_writedata,   --                                                                      .writedata
			Change_Detection_Stream_to_Mem_Translator_slave_byteenable                  => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_byteenable,  --                                                                      .byteenable
			Change_Detection_Stream_to_Mem_Translator_slave_waitrequest                 => mm_interconnect_1_change_detection_stream_to_mem_translator_slave_waitrequest  --                                                                      .waitrequest
		);

	mm_interconnect_2 : component dma_platform_mm_interconnect_2
		port map (
			System_PLL_sys_clk_clk                                                      => system_pll_sys_clk_clk,                                                                   --                                                    System_PLL_sys_clk.clk
			Change_Detection_Mem_to_Stream_Translator_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                                           -- Change_Detection_Mem_to_Stream_Translator_reset_reset_bridge_in_reset.reset
			Change_Detection_Mem_to_Stream_Translator_master_address                    => change_detection_mem_to_stream_translator_master_address,                                 --                      Change_Detection_Mem_to_Stream_Translator_master.address
			Change_Detection_Mem_to_Stream_Translator_master_waitrequest                => change_detection_mem_to_stream_translator_master_waitrequest,                             --                                                                      .waitrequest
			Change_Detection_Mem_to_Stream_Translator_master_byteenable                 => change_detection_mem_to_stream_translator_master_byteenable,                              --                                                                      .byteenable
			Change_Detection_Mem_to_Stream_Translator_master_read                       => change_detection_mem_to_stream_translator_master_read,                                    --                                                                      .read
			Change_Detection_Mem_to_Stream_Translator_master_readdata                   => change_detection_mem_to_stream_translator_master_readdata,                                --                                                                      .readdata
			Change_Detection_Mem_to_Stream_Translator_master_write                      => change_detection_mem_to_stream_translator_master_write,                                   --                                                                      .write
			Change_Detection_Mem_to_Stream_Translator_master_writedata                  => change_detection_mem_to_stream_translator_master_writedata,                               --                                                                      .writedata
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_address         => mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_address,    --           Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave.address
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_write           => mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_write,      --                                                                      .write
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_read            => mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_read,       --                                                                      .read
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_readdata        => mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_readdata,   --                                                                      .readdata
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_writedata       => mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_writedata,  --                                                                      .writedata
			Change_Detection_Mem_to_Stream_DMA_avalon_dma_control_slave_byteenable      => mm_interconnect_2_change_detection_mem_to_stream_dma_avalon_dma_control_slave_byteenable  --                                                                      .byteenable
		);

	mm_interconnect_3 : component dma_platform_mm_interconnect_3
		port map (
			System_PLL_sys_clk_clk                                                      => system_pll_sys_clk_clk,                                                                   --                                                    System_PLL_sys_clk.clk
			Change_Detection_Stream_to_Mem_Translator_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                                           -- Change_Detection_Stream_to_Mem_Translator_reset_reset_bridge_in_reset.reset
			Change_Detection_Stream_to_Mem_Translator_master_address                    => change_detection_stream_to_mem_translator_master_address,                                 --                      Change_Detection_Stream_to_Mem_Translator_master.address
			Change_Detection_Stream_to_Mem_Translator_master_waitrequest                => change_detection_stream_to_mem_translator_master_waitrequest,                             --                                                                      .waitrequest
			Change_Detection_Stream_to_Mem_Translator_master_byteenable                 => change_detection_stream_to_mem_translator_master_byteenable,                              --                                                                      .byteenable
			Change_Detection_Stream_to_Mem_Translator_master_read                       => change_detection_stream_to_mem_translator_master_read,                                    --                                                                      .read
			Change_Detection_Stream_to_Mem_Translator_master_readdata                   => change_detection_stream_to_mem_translator_master_readdata,                                --                                                                      .readdata
			Change_Detection_Stream_to_Mem_Translator_master_write                      => change_detection_stream_to_mem_translator_master_write,                                   --                                                                      .write
			Change_Detection_Stream_to_Mem_Translator_master_writedata                  => change_detection_stream_to_mem_translator_master_writedata,                               --                                                                      .writedata
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_address         => mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_address,    --           Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave.address
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_write           => mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_write,      --                                                                      .write
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_read            => mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_read,       --                                                                      .read
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_readdata        => mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_readdata,   --                                                                      .readdata
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_writedata       => mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_writedata,  --                                                                      .writedata
			Change_Detection_Stream_to_Mem_DMA_avalon_dma_control_slave_byteenable      => mm_interconnect_3_change_detection_stream_to_mem_dma_avalon_dma_control_slave_byteenable  --                                                                      .byteenable
		);

	irq_mapper : component dma_platform_irq_mapper
		port map (
			clk        => open,                    --       clk.clk
			reset      => open,                    -- clk_reset.reset
			sender_irq => arm_a9_hps_f2h_irq0_irq  --    sender.irq
		);

	irq_mapper_001 : component dma_platform_irq_mapper
		port map (
			clk        => open,                    --       clk.clk
			reset      => open,                    -- clk_reset.reset
			sender_irq => arm_a9_hps_f2h_irq1_irq  --    sender.irq
		);

	rst_controller : component dma_platform_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => arm_a9_hps_h2f_reset_reset_ports_inv, -- reset_in0.reset
			reset_in1      => system_pll_reset_source_reset,        -- reset_in1.reset
			clk            => system_pll_sys_clk_clk,               --       clk.clk
			reset_out      => rst_controller_reset_out_reset,       -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_001 : component dma_platform_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => arm_a9_hps_h2f_reset_reset_ports_inv, -- reset_in0.reset
			clk            => system_pll_sys_clk_clk,               --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,   -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_in1      => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	arm_a9_hps_h2f_reset_reset_ports_inv <= not arm_a9_hps_h2f_reset_reset;

end architecture rtl; -- of dma_platform
